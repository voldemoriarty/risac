@00000000
93 81 01 00 17 01 02 00 13 01 C1 FF 6F 00 40 1A 
13 01 01 FB 23 20 F1 02 23 26 11 04 23 24 51 04 
23 22 61 04 23 20 71 04 23 2E 81 02 23 2C 91 02 
23 2A A1 02 23 28 B1 02 23 26 C1 02 23 24 D1 02 
23 22 E1 02 23 2E 01 01 23 2C 11 01 23 2A C1 01 
23 28 D1 01 23 26 E1 01 23 24 F1 01 93 07 00 08 
73 B0 47 30 83 27 40 4B 13 07 30 06 93 87 17 00 
23 2A F0 4A 83 27 40 4B 63 8E E7 0C B7 05 00 02 
03 C5 F5 00 03 C6 05 01 83 C6 15 01 83 C7 25 01 
13 16 86 00 33 66 A6 00 93 96 06 01 B3 E6 C6 00 
93 97 87 01 B3 E7 D7 00 93 87 17 00 93 F6 F7 0F 
13 D6 87 00 03 C5 F5 00 13 87 F5 00 A3 87 D5 00 
13 76 F6 0F 93 D6 07 01 83 C5 05 01 93 F6 F6 0F 
A3 00 C7 00 03 46 27 00 23 01 D7 00 83 46 37 00 
93 D7 87 01 A3 01 F7 00 93 06 00 00 B7 07 00 03 
23 A0 D7 00 13 07 00 00 23 A2 E7 00 93 07 00 08 
73 A0 47 30 03 24 C1 03 83 20 C1 04 83 22 81 04 
03 23 41 04 83 23 01 04 83 24 81 03 03 25 41 03 
83 25 01 03 03 26 C1 02 83 26 81 02 03 27 41 02 
83 27 01 02 03 28 C1 01 83 28 81 01 03 2E 41 01 
83 2E 01 01 03 2F C1 00 83 2F 81 00 13 01 01 05 
73 00 20 30 B7 04 00 01 83 A7 44 00 93 D7 A7 00 
93 F7 17 00 E3 8C 07 F0 13 06 C0 00 93 05 C0 48 
37 05 00 01 EF 00 80 08 83 25 00 4B 37 05 00 01 
93 85 15 00 23 28 B0 4A EF 00 C0 09 13 06 20 00 
93 05 80 49 37 05 00 01 EF 00 40 06 23 2A 00 4A 
83 A7 44 00 93 E7 07 40 23 A2 F4 00 6F F0 1F ED 
13 01 01 FF 23 26 11 00 EF 00 40 1E 93 07 10 00 
63 1A F5 02 B3 86 C5 00 37 07 00 01 63 00 06 02 
83 27 47 00 93 D7 07 01 E3 8C 07 FE 83 C7 05 00 
93 85 15 00 23 00 F7 00 E3 94 B6 FE 13 05 00 00 
67 80 00 00 13 05 F0 FF 67 80 00 00 63 02 06 02 
33 87 C5 00 83 27 45 00 93 D7 07 01 E3 8C 07 FE 
83 C7 05 00 93 85 15 00 23 00 F5 00 E3 14 B7 FE 
67 80 00 00 93 07 C0 49 83 C6 07 01 83 AE 47 00 
03 AE 87 00 03 A3 C7 00 03 AF 07 00 93 D7 85 00 
13 01 01 FE 93 F7 F7 0F 23 0E D1 00 13 D6 85 01 
93 D8 47 00 93 06 01 02 93 F7 F7 00 B3 88 16 01 
13 D7 05 01 B3 86 F6 00 13 D8 C5 01 93 07 01 02 
13 76 F6 00 23 26 E1 01 23 28 D1 01 23 2A C1 01 
23 2C 61 00 13 77 F7 0F 33 88 07 01 33 86 C7 00 
93 F5 F5 0F 83 C7 C8 FE 83 CE C6 FE 03 4E C6 FE 
83 46 C8 FE 93 D8 45 00 13 08 01 02 13 56 47 00 
B3 08 18 01 33 06 C8 00 37 08 FF FF 13 08 F8 0F 
03 C3 C8 FE 93 F5 F5 00 83 48 C6 FE 13 76 F7 00 
33 F7 07 01 93 07 01 02 B3 87 B7 00 93 05 01 02 
B3 F6 06 01 33 86 C5 00 93 9E 8E 00 13 1E 8E 00 
B7 05 01 FF 93 85 F5 FF 03 C8 C7 FE 03 46 C6 FE 
B3 67 D7 01 33 E7 C6 01 B3 F7 B7 00 33 77 B7 00 
13 13 03 01 93 98 08 01 B7 06 00 01 93 86 F6 FF 
B3 E7 67 00 33 67 17 01 93 15 88 01 B3 F7 D7 00 
13 16 86 01 33 77 D7 00 B3 E7 B7 00 33 67 C7 00 
23 22 E1 00 23 24 F1 00 83 27 45 00 93 D7 07 01 
E3 8C 07 FE 93 07 00 03 23 00 F5 00 83 27 45 00 
93 D7 07 01 E3 8C 07 FE 93 07 80 07 23 00 F5 00 
13 07 41 00 93 06 C1 00 83 27 45 00 93 D7 07 01 
E3 8C 07 FE 83 47 07 00 13 07 17 00 23 00 F5 00 
E3 94 E6 FE 13 01 01 02 67 80 00 00 13 01 01 FF 
37 07 00 02 23 26 11 00 83 47 F7 00 A3 07 07 00 
83 46 07 01 23 08 07 00 83 46 17 01 A3 08 07 00 
83 46 27 01 23 09 07 00 83 27 07 00 13 07 00 40 
B7 06 00 02 13 05 00 40 63 82 E7 04 13 F6 F7 0F 
93 D5 87 00 03 C7 F6 00 93 F5 F5 0F A3 87 C6 00 
13 D6 07 01 03 C8 06 01 13 76 F6 0F 23 88 B6 00 
83 C5 16 01 93 D7 87 01 A3 88 C6 00 03 C6 26 01 
23 89 F6 00 83 A7 06 00 E3 92 A7 FC 37 07 00 02 
83 47 F7 00 A3 07 07 00 93 07 F7 00 03 47 07 01 
A3 80 07 00 03 C7 27 00 23 81 07 00 03 C7 37 00 
A3 81 07 00 93 07 00 01 73 90 57 30 93 07 00 08 
73 A0 47 30 37 05 00 01 F3 25 50 30 EF F0 9F DC 
13 06 10 00 93 05 80 49 37 05 00 01 EF F0 1F D9 
37 A6 07 00 B7 07 00 03 13 06 06 12 93 06 00 00 
23 A4 C7 00 23 A6 D7 00 6F 00 00 00 
@0000048C
49 54 53 20 41 20 54 52 41 50 3A 00 0A 00 00 00 
30 31 32 33 34 35 36 37 38 39 61 62 63 64 65 66 
00 00 00 00 
