@00000000
93 81 01 00 17 01 02 00 13 01 C1 FF 6F 00 40 00 
97 01 00 00 93 81 01 7F 17 45 00 00 13 05 05 E9 
17 46 00 00 13 06 06 EE 33 06 A6 40 93 05 00 00 
EF 00 80 2F 17 25 00 00 13 05 05 2D 63 08 05 00 
17 15 00 00 13 05 45 9B EF 20 C0 2B EF 00 40 12 
03 25 01 00 93 05 41 00 13 06 00 00 EF 30 40 42 
6F 00 C0 0D B7 47 00 00 03 C7 87 EB 63 14 07 04 
13 01 01 FF 23 24 81 00 13 84 07 00 B7 07 00 00 
23 26 11 00 93 87 07 00 63 8A 07 00 37 45 00 00 
13 05 85 EA 97 00 00 00 E7 00 00 00 93 07 10 00 
83 20 C1 00 23 0C F4 EA 03 24 81 00 13 01 01 01 
67 80 00 00 67 80 00 00 B7 07 00 00 93 87 07 00 
63 8E 07 00 B7 45 00 00 37 45 00 00 93 85 C5 EB 
13 05 85 EA 17 03 00 00 67 00 00 00 67 80 00 00 
93 07 00 00 63 94 C7 00 67 80 00 00 03 27 45 00 
13 57 07 01 E3 0C 07 FE 33 87 F5 00 03 47 07 00 
93 87 17 00 23 00 E5 00 6F F0 DF FD 93 07 10 00 
63 12 F5 02 13 01 01 FF 37 05 00 01 23 26 11 00 
EF F0 1F FC 83 20 C1 00 13 05 00 00 13 01 01 01 
67 80 00 00 13 05 F0 FF 67 80 00 00 13 01 01 FF 
93 05 00 00 23 24 81 00 23 26 11 00 13 04 05 00 
EF 00 00 42 B7 37 00 00 03 A5 07 66 83 27 C5 03 
63 84 07 00 E7 80 07 00 13 05 04 00 EF 30 00 03 
13 01 01 FF 23 24 81 00 23 20 21 01 37 04 00 00 
37 09 00 00 93 07 04 00 13 09 09 00 33 09 F9 40 
23 26 11 00 23 22 91 00 13 59 29 40 63 00 09 02 
13 04 04 00 93 04 00 00 83 27 04 00 93 84 14 00 
13 04 44 00 E7 80 07 00 E3 18 99 FE 37 04 00 00 
37 09 00 00 93 07 04 00 13 09 09 00 33 09 F9 40 
13 59 29 40 63 00 09 02 13 04 04 00 93 04 00 00 
83 27 04 00 93 84 14 00 13 04 44 00 E7 80 07 00 
E3 18 99 FE 83 20 C1 00 03 24 81 00 83 24 41 00 
03 29 01 00 13 01 01 01 67 80 00 00 B3 C7 A5 00 
93 F7 37 00 B3 08 C5 00 63 92 07 06 93 07 30 00 
63 FE C7 04 93 77 35 00 13 07 05 00 63 98 07 06 
13 F6 C8 FF 93 07 06 FE 63 6C F7 08 63 7C C7 02 
93 86 05 00 93 07 07 00 03 A8 06 00 93 87 47 00 
93 86 46 00 23 AE 07 FF E3 E8 C7 FE 93 07 F6 FF 
B3 87 E7 40 93 F7 C7 FF 93 87 47 00 33 07 F7 00 
B3 85 F5 00 63 68 17 01 67 80 00 00 13 07 05 00 
E3 7C 15 FF 83 C7 05 00 13 07 17 00 93 85 15 00 
A3 0F F7 FE E3 68 17 FF 67 80 00 00 83 C6 05 00 
13 07 17 00 93 77 37 00 A3 0F D7 FE 93 85 15 00 
E3 80 07 F8 83 C6 05 00 13 07 17 00 93 77 37 00 
A3 0F D7 FE 93 85 15 00 E3 9A 07 FC 6F F0 5F F6 
83 A6 45 00 83 A2 05 00 83 AF 85 00 03 AF C5 00 
83 AE 05 01 03 AE 45 01 03 A3 85 01 03 A8 C5 01 
23 22 D7 00 83 A6 05 02 23 20 57 00 23 24 F7 01 
23 26 E7 01 23 28 D7 01 23 2A C7 01 23 2C 67 00 
23 2E 07 01 23 20 D7 02 13 07 47 02 93 85 45 02 
E3 68 F7 FA 6F F0 9F F1 13 03 F0 00 13 07 05 00 
63 7E C3 02 93 77 F7 00 63 90 07 0A 63 92 05 08 
93 76 06 FF 13 76 F6 00 B3 86 E6 00 23 20 B7 00 
23 22 B7 00 23 24 B7 00 23 26 B7 00 13 07 07 01 
E3 66 D7 FE 63 14 06 00 67 80 00 00 B3 06 C3 40 
93 96 26 00 97 02 00 00 B3 86 56 00 67 80 C6 00 
23 07 B7 00 A3 06 B7 00 23 06 B7 00 A3 05 B7 00 
23 05 B7 00 A3 04 B7 00 23 04 B7 00 A3 03 B7 00 
23 03 B7 00 A3 02 B7 00 23 02 B7 00 A3 01 B7 00 
23 01 B7 00 A3 00 B7 00 23 00 B7 00 67 80 00 00 
93 F5 F5 0F 93 96 85 00 B3 E5 D5 00 93 96 05 01 
B3 E5 D5 00 6F F0 DF F6 93 96 27 00 97 02 00 00 
B3 86 56 00 93 82 00 00 E7 80 06 FA 93 80 02 00 
93 87 07 FF 33 07 F7 40 33 06 F6 00 E3 78 C3 F6 
6F F0 DF F3 13 01 01 FC 23 2C 81 02 13 04 05 00 
13 85 05 00 23 2A 91 02 23 2E 11 02 93 84 05 00 
EF 00 40 0C B7 37 00 00 93 87 C7 65 23 24 F1 02 
93 07 10 00 23 26 F1 02 03 27 84 03 93 07 01 02 
93 06 15 00 23 2A F1 00 93 07 20 00 23 20 91 02 
23 22 A1 02 23 2E D1 00 23 2C F1 00 83 25 84 00 
63 00 07 06 83 97 C5 00 13 97 27 01 63 42 07 02 
03 A7 45 06 B7 26 00 00 B3 E7 D7 00 B7 E6 FF FF 
93 86 F6 FF 33 77 D7 00 23 96 F5 00 23 A2 E5 06 
13 06 41 01 13 05 04 00 EF 00 80 5B 83 20 C1 03 
03 24 81 03 33 35 A0 00 33 05 A0 40 13 75 55 FF 
83 24 41 03 13 05 A5 00 13 01 01 04 67 80 00 00 
13 05 04 00 23 26 B1 00 EF 00 C0 4E 83 25 C1 00 
6F F0 5F F9 B7 47 00 00 93 05 05 00 03 A5 C7 E9 
6F F0 5F F2 93 77 35 00 13 07 05 00 63 9C 07 04 
B7 86 7F 7F 93 86 F6 F7 93 05 F0 FF 03 26 07 00 
13 07 47 00 B3 77 D6 00 B3 87 D7 00 B3 E7 C7 00 
B3 E7 D7 00 E3 84 B7 FE 83 46 C7 FF 03 46 D7 FF 
83 47 E7 FF 33 07 A7 40 63 80 06 04 63 0A 06 02 
33 35 F0 00 33 05 E5 00 13 05 E5 FF 67 80 00 00 
E3 88 06 FA 83 47 07 00 13 07 17 00 93 76 37 00 
E3 98 07 FE 33 07 A7 40 13 05 F7 FF 67 80 00 00 
13 05 D7 FF 67 80 00 00 13 05 C7 FF 67 80 00 00 
13 01 01 FD B7 37 00 00 23 2C 41 01 03 AA 07 66 
23 20 21 03 23 26 11 02 03 29 8A 14 23 24 81 02 
23 22 91 02 23 2E 31 01 23 2A 51 01 23 28 61 01 
23 26 71 01 23 24 81 01 63 00 09 04 13 0B 05 00 
93 8B 05 00 93 0A 10 00 93 09 F0 FF 83 24 49 00 
13 84 F4 FF 63 42 04 02 93 94 24 00 B3 04 99 00 
63 84 0B 04 83 A7 44 10 63 80 77 05 13 04 F4 FF 
93 84 C4 FF E3 16 34 FF 83 20 C1 02 03 24 81 02 
83 24 41 02 03 29 01 02 83 29 C1 01 03 2A 81 01 
83 2A 41 01 03 2B 01 01 83 2B C1 00 03 2C 81 00 
13 01 01 03 67 80 00 00 83 27 49 00 83 A6 44 00 
93 87 F7 FF 63 8E 87 04 23 A2 04 00 E3 88 06 FA 
83 27 89 18 33 97 8A 00 03 2C 49 00 B3 77 F7 00 
63 92 07 02 E7 80 06 00 03 27 49 00 83 27 8A 14 
63 14 87 01 E3 04 F9 F8 E3 88 07 F8 13 89 07 00 
6F F0 DF F5 83 27 C9 18 83 A5 44 08 33 77 F7 00 
63 1C 07 00 13 05 0B 00 E7 80 06 00 6F F0 DF FC 
23 22 89 00 6F F0 9F FA 13 85 05 00 E7 80 06 00 
6F F0 9F FB 13 05 00 00 67 80 00 00 B7 25 00 00 
93 85 85 37 6F 00 90 0F 13 01 01 FE 23 2E 11 00 
23 2C 81 00 23 2A 91 00 23 28 21 01 23 26 31 01 
23 24 41 01 23 22 51 01 23 20 61 01 03 24 45 00 
93 07 C0 69 23 2E F5 02 13 07 C5 2E 93 07 30 00 
23 24 E5 2E 23 22 F5 2E 23 20 05 2E 93 07 40 00 
13 09 05 00 23 26 F4 00 13 06 80 00 93 05 00 00 
23 22 04 06 23 20 04 00 23 22 04 00 23 24 04 00 
23 28 04 00 23 2A 04 00 23 2C 04 00 13 05 C4 05 
EF F0 9F C0 37 2B 00 00 83 24 89 00 B7 2A 00 00 
37 2A 00 00 B7 29 00 00 13 0B CB FD 93 8A 0A 04 
13 0A 8A 0C 93 89 09 13 B7 07 01 00 23 20 64 03 
23 22 54 03 23 24 44 03 23 26 34 03 23 2E 84 00 
93 87 97 00 23 A6 F4 00 13 06 80 00 93 05 00 00 
23 A2 04 06 23 A0 04 00 23 A2 04 00 23 A4 04 00 
23 A8 04 00 23 AA 04 00 23 AC 04 00 13 85 C4 05 
EF F0 9F B9 03 24 C9 00 B7 07 02 00 23 A0 64 03 
23 A2 54 03 23 A4 44 03 23 A6 34 03 23 AE 94 00 
93 87 27 01 23 26 F4 00 23 22 04 06 23 20 04 00 
23 22 04 00 23 24 04 00 23 28 04 00 23 2A 04 00 
23 2C 04 00 13 05 C4 05 13 06 80 00 93 05 00 00 
EF F0 9F B4 83 20 C1 01 23 20 64 03 23 22 54 03 
23 24 44 03 23 26 34 03 23 2E 84 00 03 24 81 01 
93 07 10 00 23 2C F9 02 83 24 41 01 03 29 01 01 
83 29 C1 00 03 2A 81 00 83 2A 41 00 03 2B 01 00 
13 01 01 02 67 80 00 00 13 05 00 00 67 80 00 00 
13 01 01 FF 23 22 91 00 13 06 80 06 93 84 F5 FF 
B3 84 C4 02 23 20 21 01 13 89 05 00 23 24 81 00 
23 26 11 00 93 85 44 07 EF 00 80 7F 13 04 05 00 
63 00 05 02 13 05 C5 00 23 20 04 00 23 22 24 01 
23 24 A4 00 13 86 84 06 93 05 00 00 EF F0 DF AA 
83 20 C1 00 13 05 04 00 03 24 81 00 83 24 41 00 
03 29 01 00 13 01 01 01 67 80 00 00 13 01 01 FE 
B7 37 00 00 23 28 21 01 03 A9 07 66 23 26 31 01 
23 2E 11 00 83 27 89 03 23 2C 81 00 23 2A 91 00 
93 09 05 00 63 86 07 0A 13 09 09 2E 93 04 F0 FF 
83 27 49 00 03 24 89 00 93 87 F7 FF 63 D8 07 00 
6F 00 00 08 13 04 84 06 63 8C 97 06 03 17 C4 00 
93 87 F7 FF E3 18 07 FE B7 07 FF FF 93 87 17 00 
23 22 04 06 23 20 04 00 23 22 04 00 23 24 04 00 
23 26 F4 00 23 28 04 00 23 2A 04 00 23 2C 04 00 
13 06 80 00 93 05 00 00 13 05 C4 05 EF F0 DF 9F 
23 28 04 02 23 2A 04 02 23 22 04 04 23 24 04 04 
83 20 C1 01 13 05 04 00 03 24 81 01 83 24 41 01 
03 29 01 01 83 29 C1 00 13 01 01 02 67 80 00 00 
03 24 09 00 63 0C 04 00 13 09 04 00 6F F0 5F F6 
13 05 09 00 EF F0 5F D3 6F F0 1F F5 93 05 40 00 
13 85 09 00 EF F0 DF EA 23 20 A9 00 13 04 05 00 
E3 1C 05 FC 93 07 C0 00 23 A0 F9 00 6F F0 5F FA 
B7 37 00 00 03 A5 07 66 B7 25 00 00 93 85 85 37 
6F 00 C0 5E 83 27 85 03 63 84 07 00 67 80 00 00 
6F F0 9F CE 67 80 00 00 67 80 00 00 67 80 00 00 
67 80 00 00 B7 47 00 00 03 A5 C7 E9 93 05 40 69 
6F 00 80 51 B7 47 00 00 03 A5 C7 E9 93 85 81 02 
6F 00 80 50 13 01 01 FF 23 24 81 00 B7 07 00 00 
37 04 00 00 13 04 04 00 93 87 07 00 B3 87 87 40 
23 22 91 00 23 26 11 00 93 D4 27 40 63 80 04 02 
93 87 C7 FF 33 84 87 00 83 27 04 00 93 84 F4 FF 
13 04 C4 FF E7 80 07 00 E3 98 04 FE 83 20 C1 00 
03 24 81 00 83 24 41 00 13 01 01 01 67 80 00 00 
83 27 86 00 63 8E 07 32 83 D7 C5 00 13 01 01 FD 
23 24 81 02 23 2C 41 01 23 2A 51 01 23 26 11 02 
23 22 91 02 23 20 21 03 23 2E 31 01 23 28 61 01 
23 26 71 01 23 24 81 01 23 22 91 01 23 20 A1 01 
13 F7 87 00 13 0A 06 00 93 0A 05 00 13 84 05 00 
63 06 07 08 03 A7 05 01 63 02 07 08 13 F7 27 00 
83 24 0A 00 63 0C 07 08 83 27 44 02 83 25 C4 01 
37 0B 00 80 93 09 00 00 13 09 00 00 13 4B 0B C0 
13 86 09 00 13 85 0A 00 63 02 09 04 93 06 09 00 
63 74 2B 01 93 06 0B 00 E7 80 07 00 63 58 A0 28 
83 27 8A 00 B3 89 A9 00 33 09 A9 40 33 85 A7 40 
23 24 AA 00 63 0A 05 20 83 27 44 02 83 25 C4 01 
13 86 09 00 13 85 0A 00 E3 12 09 FC 83 A9 04 00 
03 A9 44 00 93 84 84 00 6F F0 9F FA 93 05 04 00 
13 85 0A 00 EF 10 00 67 63 1C 05 3A 83 57 C4 00 
83 24 0A 00 13 F7 27 00 E3 18 07 F6 13 F7 17 00 
63 14 07 24 83 2C 84 00 03 25 04 00 37 0B 00 80 
93 4B EB FF 13 0C 00 00 13 09 00 00 13 4B FB FF 
63 0E 09 0E 13 F7 07 20 63 0C 07 24 13 8D 0C 00 
63 62 99 2F 13 F7 07 48 63 0A 07 08 83 29 44 01 
83 25 04 01 13 07 19 00 93 96 19 00 B3 86 36 01 
93 D9 F6 01 33 0D B5 40 B3 89 D9 00 93 D9 19 40 
33 07 A7 01 13 86 09 00 63 F6 E9 00 93 09 07 00 
13 06 07 00 93 F7 07 40 63 84 07 2E 93 05 06 00 
13 85 0A 00 EF 00 C0 47 93 0C 05 00 63 02 05 30 
83 25 04 01 13 06 0D 00 EF F0 4F E2 83 57 C4 00 
93 F7 F7 B7 93 E7 07 08 23 16 F4 00 33 85 AC 01 
B3 87 A9 41 23 28 94 01 23 20 A4 00 23 2A 34 01 
93 0C 09 00 23 24 F4 00 13 0D 09 00 13 06 0D 00 
93 05 0C 00 EF 00 90 4B 03 27 84 00 83 27 04 00 
93 09 09 00 B3 0C 97 41 B3 87 A7 01 23 24 94 01 
23 20 F4 00 13 09 00 00 03 26 8A 00 33 0C 3C 01 
B3 09 36 41 23 24 3A 01 63 80 09 0C 83 2C 84 00 
03 25 04 00 83 57 C4 00 E3 16 09 F0 03 AC 04 00 
03 A9 44 00 93 84 84 00 6F F0 9F EF 83 A9 44 00 
03 AC 04 00 93 84 84 00 E3 8A 09 FE 13 86 09 00 
93 05 A0 00 13 05 0C 00 EF 00 10 37 63 04 05 12 
13 05 15 00 33 0B 85 41 93 07 0B 00 93 8B 09 00 
63 F4 37 01 93 8B 07 00 03 25 04 00 83 27 04 01 
83 26 44 01 63 F8 A7 00 03 29 84 00 33 89 26 01 
63 42 79 09 63 C8 DB 1A 83 27 44 02 83 25 C4 01 
13 06 0C 00 13 85 0A 00 E7 80 07 00 13 09 05 00 
63 56 A0 08 33 0B 2B 41 13 05 10 00 63 0A 0B 16 
03 26 8A 00 33 0C 2C 01 B3 89 29 41 33 09 26 41 
23 24 2A 01 63 1A 09 08 13 05 00 00 83 20 C1 02 
03 24 81 02 83 24 41 02 03 29 01 02 83 29 C1 01 
03 2A 81 01 83 2A 41 01 03 2B 01 01 83 2B C1 00 
03 2C 81 00 83 2C 41 00 03 2D 01 00 13 01 01 03 
67 80 00 00 93 05 0C 00 13 06 09 00 EF 00 10 38 
83 27 04 00 93 05 04 00 13 85 0A 00 B3 87 27 01 
23 20 F4 00 EF 10 10 18 E3 0E 05 F6 83 17 C4 00 
93 E7 07 04 23 16 F4 00 13 05 F0 FF 6F F0 1F F9 
13 05 00 00 67 80 00 00 13 0B 00 00 13 05 00 00 
13 0C 00 00 93 09 00 00 E3 8A 09 EC E3 1E 05 EE 
13 86 09 00 93 05 A0 00 13 05 0C 00 EF 00 D0 24 
E3 10 05 EE 93 87 19 00 13 8B 07 00 6F F0 1F EE 
83 27 04 01 63 E2 A7 04 83 27 44 01 63 6E F9 02 
93 06 09 00 63 F4 2B 01 93 06 0B 00 B3 C6 F6 02 
03 27 44 02 83 25 C4 01 13 06 0C 00 13 85 0A 00 
B3 86 F6 02 E7 00 07 00 93 09 05 00 E3 58 A0 F6 
33 09 39 41 6F F0 5F E3 93 89 0C 00 63 74 99 01 
93 09 09 00 13 86 09 00 93 05 0C 00 EF 00 10 2B 
83 27 84 00 03 27 04 00 B3 87 37 41 33 07 37 01 
23 24 F4 00 23 20 E4 00 E3 94 07 FC 93 05 04 00 
13 85 0A 00 EF 10 10 0A E3 12 05 F2 33 09 39 41 
6F F0 9F DE 93 0C 09 00 13 0D 09 00 6F F0 1F DB 
93 05 04 00 13 85 0A 00 EF 10 D0 07 E3 02 05 E8 
6F F0 DF EF 13 86 0B 00 93 05 0C 00 EF 00 10 25 
83 27 84 00 03 26 04 00 13 89 0B 00 B3 87 77 41 
33 06 76 01 23 24 F4 00 23 20 C4 00 6F F0 9F E4 
13 85 0A 00 EF 00 10 35 93 0C 05 00 E3 10 05 D4 
83 25 04 01 13 85 0A 00 EF 10 50 1F 83 17 C4 00 
13 07 C0 00 23 A0 EA 00 93 F7 F7 F7 6F F0 5F EA 
13 07 C0 00 83 17 C4 00 23 A0 EA 00 6F F0 5F E9 
13 05 F0 FF 6F F0 9F E2 13 01 01 FE 23 28 21 01 
23 26 31 01 23 24 41 01 23 22 51 01 23 20 61 01 
23 2E 11 00 23 2C 81 00 23 2A 91 00 13 8B 05 00 
93 0A 05 2E 13 0A 00 00 93 09 10 00 13 09 F0 FF 
83 A4 4A 00 03 A4 8A 00 93 84 F4 FF 63 C6 04 02 
83 57 C4 00 93 84 F4 FF 63 FC F9 00 83 17 E4 00 
13 05 04 00 63 86 27 01 E7 00 0B 00 33 6A AA 00 
13 04 84 06 E3 9E 24 FD 83 AA 0A 00 E3 92 0A FC 
83 20 C1 01 03 24 81 01 83 24 41 01 03 29 01 01 
83 29 C1 00 83 2A 41 00 03 2B 01 00 13 05 0A 00 
03 2A 81 00 13 01 01 02 67 80 00 00 13 01 01 FD 
23 20 21 03 23 2E 31 01 23 2C 41 01 23 2A 51 01 
23 28 61 01 23 26 71 01 23 26 11 02 23 24 81 02 
23 22 91 02 93 0A 05 00 93 8B 05 00 13 0B 05 2E 
13 0A 00 00 93 09 10 00 13 09 F0 FF 83 24 4B 00 
03 24 8B 00 93 84 F4 FF 63 C8 04 02 83 57 C4 00 
93 84 F4 FF 63 FE F9 00 83 17 E4 00 93 05 04 00 
13 85 0A 00 63 86 27 01 E7 80 0B 00 33 6A AA 00 
13 04 84 06 E3 9C 24 FD 03 2B 0B 00 E3 10 0B FC 
83 20 C1 02 03 24 81 02 83 24 41 02 03 29 01 02 
83 29 C1 01 83 2A 41 01 03 2B 01 01 83 2B C1 00 
13 05 0A 00 03 2A 81 01 13 01 01 03 67 80 00 00 
13 01 01 FD 23 2E 31 01 23 26 11 02 23 24 81 02 
23 22 91 02 23 20 21 03 23 2C 41 01 23 2A 51 01 
23 28 61 01 23 26 71 01 23 24 81 01 23 22 91 01 
93 87 B5 00 13 07 60 01 93 09 05 00 63 66 F7 06 
93 07 00 01 63 E6 B7 1E EF 00 50 16 93 04 00 01 
13 06 20 00 93 07 80 01 37 49 00 00 13 09 09 A9 
B3 07 F9 00 03 A4 47 00 13 87 87 FF 63 0A E4 20 
83 27 44 00 83 26 C4 00 03 26 84 00 93 F7 C7 FF 
B3 07 F4 00 03 A7 47 00 23 26 D6 00 23 A4 C6 00 
13 67 17 00 13 85 09 00 23 A2 E7 00 EF 00 50 11 
13 05 84 00 6F 00 80 19 93 F4 87 FF 63 C2 07 18 
63 E0 B4 18 EF 00 90 0F 93 07 70 1F 63 F6 97 46 
93 D7 94 00 63 86 07 1A 13 07 40 00 63 6C F7 3C 
93 D7 64 00 13 86 97 03 13 85 87 03 93 16 36 00 
37 49 00 00 13 09 09 A9 B3 06 D9 00 03 A4 46 00 
93 86 86 FF 63 86 86 02 93 05 F0 00 6F 00 00 01 
63 5C 07 32 03 24 C4 00 63 8C 86 00 83 27 44 00 
93 F7 C7 FF 33 87 97 40 E3 D4 E5 FE 13 06 05 00 
03 24 09 01 93 08 89 00 63 08 14 17 03 25 44 00 
93 06 F0 00 13 75 C5 FF B3 07 95 40 63 CC F6 40 
23 2A 19 01 23 28 19 01 63 D6 07 3E 93 07 F0 1F 
63 EA A7 2E 93 77 85 FF 93 87 87 00 83 25 49 00 
B3 07 F9 00 83 A6 07 00 13 55 55 00 13 07 10 00 
33 17 A7 00 33 67 B7 00 93 85 87 FF 23 26 B4 00 
23 24 D4 00 23 22 E9 00 23 A0 87 00 23 A6 86 00 
93 57 26 40 93 05 10 00 B3 95 F5 00 63 68 B7 10 
B3 F7 E5 00 63 94 07 02 93 95 15 00 13 76 C6 FF 
B3 F7 E5 00 13 06 46 00 63 9A 07 00 93 95 15 00 
B3 F7 E5 00 13 06 46 00 E3 8A 07 FE 13 08 F0 00 
13 13 36 00 33 03 69 00 13 05 03 00 83 27 C5 00 
13 0E 06 00 63 02 F5 2E 03 A7 47 00 13 84 07 00 
83 A7 C7 00 13 77 C7 FF B3 06 97 40 63 42 D8 2E 
E3 C2 06 FE 33 07 E4 00 83 26 47 00 03 26 84 00 
13 85 09 00 93 E6 16 00 23 22 D7 00 23 26 F6 00 
23 A4 C7 00 EF 00 C0 78 13 05 84 00 6F 00 00 01 
93 07 C0 00 23 A0 F9 00 13 05 00 00 83 20 C1 02 
03 24 81 02 83 24 41 02 03 29 01 02 83 29 C1 01 
03 2A 81 01 83 2A 41 01 03 2B 01 01 83 2B C1 00 
03 2C 81 00 83 2C 41 00 13 01 01 03 67 80 00 00 
93 06 00 20 13 06 00 04 13 05 F0 03 6F F0 5F E6 
03 A4 C7 00 13 06 26 00 E3 94 87 DE 03 24 09 01 
93 08 89 00 E3 1C 14 E9 03 27 49 00 93 57 26 40 
93 05 10 00 B3 95 F5 00 E3 7C B7 EE 03 24 89 00 
83 2A 44 00 13 FB CA FF 63 68 9B 00 B3 07 9B 40 
13 07 F0 00 63 46 F7 14 B7 47 00 00 B7 4C 00 00 
83 AA 87 F0 03 A7 0C EA 93 07 F0 FF 33 0A 64 01 
B3 8A 54 01 63 0A F7 34 B7 17 00 00 93 87 F7 00 
B3 8A FA 00 B7 F7 FF FF B3 FA FA 00 93 85 0A 00 
13 85 09 00 EF 00 90 42 93 07 F0 FF 93 0B 05 00 
63 0C F5 28 63 68 45 29 37 4C 00 00 13 0C 4C ED 
83 25 0C 00 B3 85 BA 00 23 20 BC 00 93 87 05 00 
63 04 AA 3A 83 A6 0C EA 13 07 F0 FF 63 8C E6 3A 
33 8A 4B 41 B3 07 FA 00 23 20 FC 00 93 FC 7B 00 
63 86 0C 30 B7 17 00 00 B3 8B 9B 41 93 85 87 00 
93 8B 8B 00 B3 85 95 41 B3 8A 5B 01 93 87 F7 FF 
B3 85 55 41 33 FA F5 00 93 05 0A 00 13 85 09 00 
EF 00 D0 3A 93 07 F0 FF 63 00 F5 3C 33 05 75 41 
B3 0A 45 01 83 25 0C 00 23 24 79 01 93 EA 1A 00 
B3 05 BA 00 23 20 BC 00 23 A2 5B 01 63 08 24 35 
93 06 F0 00 63 F8 66 35 03 27 44 00 93 07 4B FF 
93 F7 87 FF 13 77 17 00 33 67 F7 00 23 22 E4 00 
13 06 50 00 33 07 F4 00 23 22 C7 00 23 24 C7 00 
63 EE F6 36 83 AA 4B 00 13 84 0B 00 B7 47 00 00 
03 A7 47 F0 63 74 B7 00 23 A2 B7 F0 B7 47 00 00 
03 A7 07 F0 63 76 B7 1A 23 A0 B7 F0 6F 00 40 1A 
13 E7 14 00 23 22 E4 00 B3 04 94 00 23 24 99 00 
93 E7 17 00 13 85 09 00 23 A2 F4 00 EF 00 40 58 
13 05 84 00 6F F0 9F E0 83 26 C4 00 03 26 84 00 
6F F0 1F C4 93 57 95 00 13 07 40 00 63 72 F7 14 
13 07 40 01 63 6A F7 22 93 86 C7 05 93 85 B7 05 
93 96 36 00 B3 06 D9 00 83 A7 06 00 93 86 86 FF 
63 88 F6 1C 03 A7 47 00 13 77 C7 FF 63 76 E5 00 
83 A7 87 00 E3 98 F6 FE 83 A6 C7 00 03 27 49 00 
23 26 D4 00 23 24 F4 00 23 A4 86 00 23 A6 87 00 
6F F0 1F CF 13 07 40 01 63 76 F7 12 13 07 40 05 
63 6A F7 1E 93 D7 C4 00 13 86 F7 06 13 85 E7 06 
93 16 36 00 6F F0 DF C1 13 0E 1E 00 93 77 3E 00 
13 05 85 00 63 8E 07 10 83 27 C5 00 6F F0 9F D0 
03 26 84 00 93 E5 14 00 23 22 B4 00 23 26 F6 00 
23 A4 C7 00 B3 04 94 00 23 2A 99 00 23 28 99 00 
93 E7 16 00 23 A6 14 01 23 A4 14 01 23 A2 F4 00 
33 07 E4 00 13 85 09 00 23 20 D7 00 EF 00 40 49 
13 05 84 00 6F F0 9F D1 13 D6 34 00 93 87 84 00 
6F F0 9F B2 33 07 A4 00 83 27 47 00 13 85 09 00 
93 E7 17 00 23 22 F7 00 EF 00 80 46 13 05 84 00 
6F F0 DF CE 13 E7 14 00 23 22 E4 00 B3 04 94 00 
23 2A 99 00 23 28 99 00 13 E7 17 00 23 A6 14 01 
23 A4 14 01 23 A2 E4 00 33 05 A4 00 23 20 F5 00 
13 85 09 00 EF 00 C0 42 13 05 84 00 6F F0 1F CB 
93 57 65 00 93 86 97 03 93 85 87 03 93 96 36 00 
6F F0 5F EC 63 0E 24 11 03 24 89 00 83 2A 44 00 
93 FA CA FF B3 87 9A 40 63 E6 9A 00 13 07 F0 00 
E3 48 F7 E4 13 85 09 00 EF 00 80 3E 13 05 00 00 
6F F0 DF C6 13 86 C7 05 13 85 B7 05 93 16 36 00 
6F F0 1F B0 83 27 83 00 13 06 F6 FF 63 92 67 1C 
93 77 36 00 13 03 83 FF E3 96 07 FE 03 27 49 00 
93 C7 F5 FF B3 F7 E7 00 23 22 F9 00 93 95 15 00 
E3 EE B7 C8 E3 8C 05 C8 33 F7 F5 00 63 1A 07 00 
93 95 15 00 33 F7 F5 00 13 0E 4E 00 E3 0A 07 FE 
13 06 0E 00 6F F0 DF B9 93 8A 0A 01 6F F0 1F CC 
03 25 49 00 93 D5 25 40 13 07 10 00 33 17 B7 00 
33 67 A7 00 23 22 E9 00 6F F0 9F E3 B3 85 5B 01 
B3 05 B0 40 93 95 45 01 13 DA 45 01 93 05 0A 00 
13 85 09 00 EF 00 90 0B 93 07 F0 FF E3 18 F5 D0 
13 0A 00 00 6F F0 1F D1 13 07 40 05 63 62 F7 08 
93 57 C5 00 93 86 F7 06 93 85 E7 06 93 96 36 00 
6F F0 5F DC 13 07 40 15 63 62 F7 08 93 D7 F4 00 
13 86 87 07 13 85 77 07 93 16 36 00 6F F0 5F A2 
37 4C 00 00 13 0C 4C ED 83 27 0C 00 B3 87 FA 00 
23 20 FC 00 6F F0 1F C6 13 17 4A 01 E3 1C 07 C4 
03 24 89 00 B3 0A 5B 01 93 EA 1A 00 23 22 54 01 
6F F0 DF CF 23 A0 7C EB 6F F0 5F C5 13 84 0B 00 
6F F0 DF CE 93 07 10 00 23 A2 FB 00 6F F0 9F EB 
13 07 40 15 63 62 F7 06 93 57 F5 00 93 86 87 07 
93 85 77 07 93 96 36 00 6F F0 DF D3 13 07 40 55 
63 62 F7 06 93 D7 24 01 13 86 D7 07 13 85 C7 07 
93 16 36 00 6F F0 DF 99 93 8C 8C FF B3 8A 9A 01 
B3 8A 7A 41 13 0A 00 00 6F F0 DF C3 93 05 84 00 
13 85 09 00 EF 10 80 10 03 24 89 00 83 25 0C 00 
83 2A 44 00 6F F0 9F C7 13 07 40 55 63 64 F7 02 
93 57 25 01 93 86 D7 07 93 85 C7 07 93 96 36 00 
6F F0 5F CD 93 06 80 3F 13 06 F0 07 13 05 E0 07 
6F F0 1F 94 93 06 80 3F 93 05 E0 07 6F F0 9F CB 
83 27 49 00 6F F0 9F E5 93 77 35 00 93 F6 F5 0F 
63 8A 07 02 93 07 F6 FF 63 0E 06 02 13 06 F0 FF 
6F 00 80 01 13 05 15 00 13 77 35 00 63 0E 07 00 
93 87 F7 FF 63 80 C7 02 03 47 05 00 E3 14 D7 FE 
67 80 00 00 93 07 06 00 13 07 30 00 63 66 F7 02 
63 96 07 00 13 05 00 00 67 80 00 00 B3 07 F5 00 
6F 00 C0 00 13 05 15 00 E3 86 A7 FE 03 47 05 00 
E3 1A D7 FE 67 80 00 00 37 07 01 00 93 98 85 00 
13 07 F7 FF B3 F8 E8 00 93 F5 F5 0F B3 E5 B8 00 
93 98 05 01 B3 E8 B8 00 37 08 FF FE B7 85 80 80 
13 08 F8 EF 93 85 05 08 13 03 30 00 03 27 05 00 
33 C7 E8 00 33 06 07 01 13 47 F7 FF 33 77 E6 00 
33 77 B7 00 E3 1C 07 F8 93 87 C7 FF 13 05 45 00 
E3 6E F3 FC E3 94 07 F8 6F F0 DF F7 63 F6 A5 02 
B3 87 C5 00 63 72 F5 02 33 07 C5 00 63 0A 06 0E 
83 C6 F7 FF 93 87 F7 FF 13 07 F7 FF 23 00 D7 00 
E3 98 F5 FE 67 80 00 00 93 07 F0 00 63 E8 C7 02 
93 07 05 00 93 06 F6 FF 63 0C 06 0C 93 86 16 00 
B3 86 D7 00 03 C7 05 00 93 87 17 00 93 85 15 00 
A3 8F E7 FE E3 98 D7 FE 67 80 00 00 B3 E7 A5 00 
93 F7 37 00 63 90 07 0A 93 08 06 FF 93 F8 08 FF 
93 88 08 01 33 08 15 01 13 87 05 00 93 07 05 00 
83 26 07 00 13 07 07 01 93 87 07 01 23 A8 D7 FE 
83 26 47 FF 23 AA D7 FE 83 26 87 FF 23 AC D7 FE 
83 26 C7 FF 23 AE D7 FE E3 1C F8 FC 13 77 C6 00 
B3 85 15 01 13 78 F6 00 63 0E 07 04 13 87 05 00 
93 88 07 00 13 0E 30 00 03 23 07 00 13 07 47 00 
B3 06 E8 40 23 A0 68 00 B3 86 D5 00 93 88 48 00 
E3 64 DE FE 13 07 C8 FF 13 77 C7 FF 13 07 47 00 
13 76 36 00 B3 87 E7 00 B3 85 E5 00 6F F0 9F F3 
67 80 00 00 93 06 F6 FF 93 07 05 00 6F F0 1F F3 
67 80 00 00 13 06 08 00 6F F0 DF F1 67 80 00 00 
67 80 00 00 13 01 01 FD 23 20 21 03 23 26 11 02 
23 24 81 02 23 22 91 02 23 2E 31 01 23 2C 41 01 
23 2A 51 01 23 28 61 01 23 26 71 01 23 24 81 01 
13 09 06 00 63 84 05 22 13 84 05 00 93 09 05 00 
EF F0 DF FB 93 04 B9 00 93 07 60 01 63 FE 97 0E 
93 F4 84 FF 13 87 04 00 63 CE 04 0E 63 EC 24 0F 
83 27 C4 FF 93 0A 84 FF 13 FA C7 FF 33 8B 4A 01 
63 5C EA 18 B7 46 00 00 93 8B 06 A9 03 A6 8B 00 
83 26 4B 00 63 0E 66 23 13 F6 E6 FF 33 06 CB 00 
03 26 46 00 13 76 16 00 63 14 06 1A 93 F6 C6 FF 
33 06 DA 00 63 5E E6 32 93 F7 17 00 63 94 07 02 
03 2C 84 FF 33 8C 8A 41 83 27 4C 00 93 F7 C7 FF 
B3 86 D7 00 B3 8B 46 01 63 DA EB 34 B3 0B FA 00 
63 D2 EB 0C 93 05 09 00 13 85 09 00 EF F0 4F D7 
13 09 05 00 63 0C 05 04 83 27 C4 FF 13 07 85 FF 
93 F7 E7 FF B3 87 FA 00 63 82 E7 30 13 06 CA FF 
93 07 40 02 63 E6 C7 30 13 07 30 01 83 26 04 00 
63 6C C7 26 93 07 05 00 13 07 04 00 23 A0 D7 00 
83 26 47 00 23 A2 D7 00 03 27 87 00 23 A4 E7 00 
93 05 04 00 13 85 09 00 EF 00 50 58 13 85 09 00 
EF F0 1F EC 6F 00 C0 01 93 04 00 01 13 07 00 01 
E3 F8 24 F1 93 07 C0 00 23 A0 F9 00 13 09 00 00 
83 20 C1 02 03 24 81 02 83 24 41 02 83 29 C1 01 
03 2A 81 01 83 2A 41 01 03 2B 01 01 83 2B C1 00 
03 2C 81 00 13 05 09 00 03 29 01 02 13 01 01 03 
67 80 00 00 83 27 CC 00 03 27 8C 00 13 06 CA FF 
93 06 40 02 23 26 F7 00 23 A4 E7 00 13 09 8C 00 
33 0B 7C 01 63 E4 C6 2E 93 05 30 01 03 27 04 00 
93 07 09 00 63 F2 C5 02 23 24 EC 00 03 27 44 00 
93 07 B0 01 23 26 EC 00 63 E2 C7 30 03 27 84 00 
93 07 0C 01 13 04 84 00 23 A0 E7 00 03 27 44 00 
13 8A 0B 00 93 0A 0C 00 23 A2 E7 00 03 27 84 00 
13 04 09 00 23 A4 E7 00 83 A7 4A 00 33 07 9A 40 
93 06 F0 00 93 F7 17 00 63 EC E6 06 B3 67 FA 00 
23 A2 FA 00 83 27 4B 00 93 E7 17 00 23 22 FB 00 
13 85 09 00 EF F0 DF DC 13 09 04 00 6F F0 5F F2 
93 F7 17 00 E3 98 07 E8 03 2C 84 FF 33 8C 8A 41 
83 27 4C 00 93 F7 C7 FF 6F F0 5F E7 03 24 81 02 
83 20 C1 02 83 24 41 02 03 29 01 02 83 29 C1 01 
03 2A 81 01 83 2A 41 01 03 2B 01 01 83 2B C1 00 
03 2C 81 00 93 05 06 00 13 01 01 03 6F F0 4F BC 
B3 E7 97 00 23 A2 FA 00 B3 85 9A 00 13 67 17 00 
23 A2 E5 00 83 27 4B 00 93 85 85 00 13 85 09 00 
93 E7 17 00 23 22 FB 00 EF 00 50 40 6F F0 5F F7 
93 F6 C6 FF 33 06 DA 00 93 85 04 01 63 50 B6 0E 
93 F7 17 00 E3 90 07 E0 03 2C 84 FF 33 8C 8A 41 
83 27 4C 00 93 F7 C7 FF B3 86 D7 00 33 8B 46 01 
E3 4E BB DC 83 27 CC 00 03 27 8C 00 13 06 CA FF 
93 06 40 02 23 26 F7 00 23 A4 E7 00 13 09 8C 00 
63 EE C6 20 93 05 30 01 03 27 04 00 93 07 09 00 
63 F2 C5 02 23 24 EC 00 03 27 44 00 93 07 B0 01 
23 26 EC 00 63 E4 C7 20 03 27 84 00 93 07 0C 01 
13 04 84 00 23 A0 E7 00 03 27 44 00 23 A2 E7 00 
03 27 84 00 23 A4 E7 00 33 07 9C 00 B3 07 9B 40 
23 A4 EB 00 93 E7 17 00 23 22 F7 00 83 27 4C 00 
13 85 09 00 93 F7 17 00 B3 E4 97 00 23 22 9C 00 
EF F0 1F C8 6F F0 DF DD 23 20 D5 00 83 26 44 00 
13 07 B0 01 23 22 D5 00 63 60 C7 12 83 26 84 00 
13 07 84 00 93 07 85 00 6F F0 5F D7 B3 8A 9A 00 
B3 07 96 40 23 A4 5B 01 93 E7 17 00 23 A2 FA 00 
83 27 C4 FF 13 85 09 00 13 09 04 00 93 F7 17 00 
B3 E4 97 00 23 2E 94 FE EF F0 9F C2 6F F0 5F D8 
83 27 CB 00 03 27 8B 00 13 0A 06 00 33 8B CA 00 
23 26 F7 00 23 A4 E7 00 6F F0 1F E1 83 27 C5 FF 
93 F7 C7 FF 33 0A FA 00 33 8B 4A 01 6F F0 DF DF 
93 05 04 00 EF F0 9F AC 6F F0 9F D1 83 27 CB 00 
03 27 8B 00 13 06 CA FF 93 06 40 02 23 26 F7 00 
23 A4 E7 00 03 27 8C 00 83 27 CC 00 13 09 8C 00 
33 0B 7C 01 23 26 F7 00 23 A4 E7 00 63 E8 C6 04 
93 06 30 01 03 27 04 00 93 07 09 00 E3 F6 C6 D8 
23 24 EC 00 03 27 44 00 93 07 B0 01 23 26 EC 00 
03 27 84 00 E3 F6 C7 D6 23 28 EC 00 03 27 C4 00 
93 07 40 02 23 2A EC 00 03 27 04 01 63 04 F6 06 
93 07 8C 01 13 04 04 01 6F F0 1F D5 93 05 04 00 
13 05 09 00 EF F0 9F A3 13 04 09 00 13 8A 0B 00 
93 0A 0C 00 6F F0 5F D5 03 27 84 00 23 24 E5 00 
03 27 C4 00 23 26 E5 00 83 26 04 01 63 02 F6 04 
13 07 04 01 93 07 05 01 6F F0 5F C4 83 27 84 00 
23 28 FC 00 83 27 C4 00 23 2A FC 00 03 27 04 01 
E3 10 D6 FA 23 2C EC 00 03 27 44 01 93 07 0C 02 
13 04 84 01 23 2E EC 00 03 27 04 00 6F F0 DF CD 
23 28 D5 00 83 26 44 01 13 07 84 01 93 07 85 01 
23 2A D5 00 83 26 84 01 6F F0 5F BF 93 05 04 00 
13 05 09 00 EF F0 9F 9A 6F F0 1F E2 83 27 84 00 
23 28 FC 00 83 27 C4 00 23 2A FC 00 03 27 04 01 
63 08 D6 00 93 07 8C 01 13 04 04 01 6F F0 9F DE 
23 2C EC 00 03 27 44 01 93 07 0C 02 13 04 84 01 
23 2E EC 00 03 27 04 00 6F F0 DF DC 13 01 01 FF 
23 24 81 00 23 22 91 00 13 04 05 00 B7 44 00 00 
13 85 05 00 23 26 11 00 23 AE 04 EE EF 10 40 39 
93 07 F0 FF 63 0C F5 00 83 20 C1 00 03 24 81 00 
83 24 41 00 13 01 01 01 67 80 00 00 83 A7 C4 EF 
E3 84 07 FE 83 20 C1 00 23 20 F4 00 03 24 81 00 
83 24 41 00 13 01 01 01 67 80 00 00 13 01 01 FF 
23 24 81 00 13 84 05 00 83 95 E5 00 23 26 11 00 
EF 00 90 63 63 40 05 02 83 27 04 05 83 20 C1 00 
B3 87 A7 00 23 28 F4 04 03 24 81 00 13 01 01 01 
67 80 00 00 83 57 C4 00 37 F7 FF FF 13 07 F7 FF 
B3 F7 E7 00 83 20 C1 00 23 16 F4 00 03 24 81 00 
13 01 01 01 67 80 00 00 13 05 00 00 67 80 00 00 
83 97 C5 00 13 01 01 FE 23 2C 81 00 23 2A 91 00 
23 28 21 01 23 26 31 01 23 2E 11 00 13 F7 07 10 
13 84 05 00 93 04 05 00 83 95 E5 00 13 09 06 00 
93 89 06 00 63 1E 07 02 37 F7 FF FF 13 07 F7 FF 
B3 F7 E7 00 23 16 F4 00 03 24 81 01 83 20 C1 01 
93 86 09 00 13 06 09 00 83 29 C1 00 03 29 01 01 
13 85 04 00 83 24 41 01 13 01 01 02 6F 00 C0 08 
93 06 20 00 13 06 00 00 EF 00 90 31 83 17 C4 00 
83 15 E4 00 6F F0 5F FB 13 01 01 FF 23 24 81 00 
13 84 05 00 83 95 E5 00 23 26 11 00 EF 00 50 2F 
93 07 F0 FF 63 04 F5 02 83 57 C4 00 37 17 00 00 
83 20 C1 00 B3 E7 E7 00 23 28 A4 04 23 16 F4 00 
03 24 81 00 13 01 01 01 67 80 00 00 83 57 C4 00 
37 F7 FF FF 13 07 F7 FF B3 F7 E7 00 83 20 C1 00 
23 16 F4 00 03 24 81 00 13 01 01 01 67 80 00 00 
83 95 E5 00 6F 00 40 1E 13 01 01 FF 13 87 05 00 
23 24 81 00 23 22 91 00 93 05 06 00 13 04 05 00 
B7 44 00 00 13 86 06 00 13 05 07 00 23 26 11 00 
23 AE 04 EE EF D0 9F FA 93 07 F0 FF 63 0C F5 00 
83 20 C1 00 03 24 81 00 83 24 41 00 13 01 01 01 
67 80 00 00 83 A7 C4 EF E3 84 07 FE 83 20 C1 00 
23 20 F4 00 03 24 81 00 83 24 41 00 13 01 01 01 
67 80 00 00 B7 47 00 00 83 A7 C7 E9 13 01 01 FF 
23 24 81 00 23 22 91 00 23 26 11 00 93 04 05 00 
13 84 05 00 63 86 07 00 03 A7 87 03 63 00 07 0E 
03 17 C4 00 93 17 07 01 93 76 87 00 93 D7 07 01 
63 80 06 04 83 26 04 01 63 80 06 06 13 F6 17 00 
63 04 06 08 03 26 44 01 23 24 04 00 13 05 00 00 
33 06 C0 40 23 2C C4 00 63 86 06 08 83 20 C1 00 
03 24 81 00 83 24 41 00 13 01 01 01 67 80 00 00 
93 F6 07 01 63 84 06 0C 93 F7 47 00 63 96 07 08 
83 26 04 01 13 67 87 00 93 17 07 01 23 16 E4 00 
93 D7 07 01 E3 94 06 FA 13 F6 07 28 93 05 00 20 
E3 0E B6 F8 93 05 04 00 13 85 04 00 EF 00 10 2B 
03 17 C4 00 83 26 04 01 93 17 07 01 93 D7 07 01 
13 F6 17 00 E3 10 06 F8 13 F6 27 00 93 05 00 00 
63 14 06 00 83 25 44 01 23 24 B4 00 13 05 00 00 
E3 9E 06 F6 93 F7 07 08 E3 8A 07 F6 13 67 07 04 
23 16 E4 00 13 05 F0 FF 6F F0 5F F6 13 85 07 00 
EF E0 4F F0 6F F0 DF F1 83 25 04 03 63 8E 05 00 
93 07 04 04 63 88 F5 00 13 85 04 00 EF 00 00 5F 
03 17 C4 00 23 28 04 02 83 26 04 01 13 77 B7 FD 
23 22 04 00 23 20 D4 00 6F F0 DF F4 93 07 90 00 
23 A0 F4 00 13 67 07 04 23 16 E4 00 13 05 F0 FF 
6F F0 DF F0 93 05 05 00 93 06 00 00 13 06 00 00 
13 05 00 00 6F 00 D0 4C 13 01 01 FF 23 24 81 00 
23 22 91 00 13 04 05 00 B7 44 00 00 13 85 05 00 
23 26 11 00 23 AE 04 EE EF 00 D0 60 93 07 F0 FF 
63 0C F5 00 83 20 C1 00 03 24 81 00 83 24 41 00 
13 01 01 01 67 80 00 00 83 A7 C4 EF E3 84 07 FE 
83 20 C1 00 23 20 F4 00 03 24 81 00 83 24 41 00 
13 01 01 01 67 80 00 00 13 01 01 FF 23 26 11 00 
23 24 81 00 23 22 91 00 23 20 21 01 63 80 05 02 
13 84 05 00 93 04 05 00 63 06 05 00 83 27 85 03 
63 8C 07 0A 83 17 C4 00 63 92 07 02 83 20 C1 00 
03 24 81 00 13 09 00 00 83 24 41 00 13 05 09 00 
03 29 01 00 13 01 01 01 67 80 00 00 93 05 04 00 
13 85 04 00 EF 00 40 0C 83 27 C4 02 13 09 05 00 
63 8A 07 00 83 25 C4 01 13 85 04 00 E7 80 07 00 
63 4C 05 06 83 57 C4 00 93 F7 07 08 63 9E 07 06 
83 25 04 03 63 8C 05 00 93 07 04 04 63 86 F5 00 
13 85 04 00 EF 00 80 4A 23 28 04 02 83 25 44 04 
63 88 05 00 13 85 04 00 EF 00 40 49 23 22 04 04 
EF E0 4F D9 23 16 04 00 EF E0 0F D9 83 20 C1 00 
03 24 81 00 83 24 41 00 13 05 09 00 03 29 01 00 
13 01 01 01 67 80 00 00 EF E0 CF D5 83 17 C4 00 
E3 86 07 F4 6F F0 9F F6 83 57 C4 00 13 09 F0 FF 
93 F7 07 08 E3 86 07 F8 83 25 04 01 13 85 04 00 
EF 00 C0 43 6F F0 DF F7 B7 47 00 00 93 05 05 00 
03 A5 C7 E9 6F F0 5F EE 83 97 C5 00 13 01 01 FE 
23 2C 81 00 23 26 31 01 23 2E 11 00 23 2A 91 00 
23 28 21 01 93 F6 87 00 13 84 05 00 93 09 05 00 
63 9A 06 10 37 17 00 00 13 07 07 80 83 A6 45 00 
B3 E7 E7 00 23 96 F5 00 63 54 D0 18 03 27 84 02 
63 0A 07 0C 83 A4 09 00 93 96 07 01 23 A0 09 00 
13 96 37 01 83 25 C4 01 93 D6 06 01 63 48 06 16 
93 06 10 00 13 06 00 00 13 85 09 00 E7 00 07 00 
93 07 F0 FF 63 0C F5 18 83 56 C4 00 03 27 84 02 
83 25 C4 01 93 F6 46 00 63 8E 06 00 83 26 44 00 
83 27 04 03 33 05 D5 40 63 86 07 00 83 27 C4 03 
33 05 F5 40 13 06 05 00 93 06 00 00 13 85 09 00 
E7 00 07 00 93 07 F0 FF 63 1E F5 10 03 A7 09 00 
83 17 C4 00 63 08 07 16 93 06 D0 01 63 06 D7 00 
93 06 60 01 63 14 D7 0C 83 26 04 01 37 F7 FF FF 
13 07 F7 7F B3 F7 E7 00 23 16 F4 00 23 22 04 00 
23 20 D4 00 83 25 04 03 23 A0 99 00 63 8C 05 00 
93 07 04 04 63 86 F5 00 13 85 09 00 EF 00 00 31 
23 28 04 02 13 05 00 00 83 20 C1 01 03 24 81 01 
83 24 41 01 03 29 01 01 83 29 C1 00 13 01 01 02 
67 80 00 00 03 A9 05 01 E3 0E 09 FC 83 A4 05 00 
13 97 07 01 13 57 07 01 13 77 37 00 23 A0 25 01 
B3 84 24 41 93 07 00 00 63 14 07 00 83 A7 45 01 
23 24 F4 00 63 48 90 00 6F F0 DF FA 33 09 A9 00 
E3 52 90 FA 83 27 44 02 83 25 C4 01 93 86 04 00 
13 06 09 00 13 85 09 00 E7 80 07 00 B3 84 A4 40 
E3 4E A0 FC 83 57 C4 00 13 05 F0 FF 93 E7 07 04 
83 20 C1 01 23 16 F4 00 03 24 81 01 83 24 41 01 
03 29 01 01 83 29 C1 00 13 01 01 02 67 80 00 00 
03 A7 C5 03 E3 4C E0 E6 6F F0 DF F4 03 25 04 05 
6F F0 5F EB 83 57 C4 00 37 F7 FF FF 13 07 F7 7F 
B3 F7 E7 00 83 26 04 01 93 97 07 01 93 D7 07 41 
23 16 F4 00 23 22 04 00 23 20 D4 00 13 97 37 01 
E3 5A 07 EE 23 28 A4 04 6F F0 DF EE 83 A7 09 00 
E3 84 07 E6 13 07 D0 01 63 88 E7 02 13 07 60 01 
63 84 E7 02 83 57 C4 00 93 E7 07 04 23 16 F4 00 
6F F0 9F EE 37 F7 FF FF 13 07 F7 7F 83 26 04 01 
B3 F7 E7 00 6F F0 DF FA 23 A0 99 00 13 05 00 00 
6F F0 9F EC 13 01 01 FE 23 2C 81 00 23 2E 11 00 
13 04 05 00 63 06 05 00 83 27 85 03 63 80 07 02 
83 97 C5 00 63 96 07 02 83 20 C1 01 03 24 81 01 
13 05 00 00 13 01 01 02 67 80 00 00 23 26 B1 00 
EF E0 4F A8 83 25 C1 00 83 97 C5 00 E3 8E 07 FC 
13 05 04 00 03 24 81 01 83 20 C1 01 13 01 01 02 
6F F0 9F D4 93 05 05 00 63 08 05 00 B7 47 00 00 
03 A5 C7 E9 6F F0 1F F9 B7 37 00 00 03 A5 07 66 
B7 25 00 00 93 85 45 6F 6F E0 5F 82 13 01 01 FE 
23 26 31 01 B7 49 00 00 23 2C 81 00 23 2A 91 00 
23 28 21 01 23 24 41 01 23 2E 11 00 13 8A 05 00 
13 09 05 00 93 89 09 A9 EF F0 4F A5 03 A7 89 00 
B7 17 00 00 13 84 F7 FE 83 24 47 00 33 04 44 41 
93 F4 C4 FF 33 04 94 00 13 54 C4 00 13 04 F4 FF 
13 14 C4 00 63 4E F4 00 93 05 00 00 13 05 09 00 
EF F0 CF F9 83 A7 89 00 B3 87 97 00 63 08 F5 02 
13 05 09 00 EF F0 CF A0 83 20 C1 01 03 24 81 01 
83 24 41 01 03 29 01 01 83 29 C1 00 03 2A 81 00 
13 05 00 00 13 01 01 02 67 80 00 00 B3 05 80 40 
13 05 09 00 EF F0 8F F5 93 07 F0 FF 63 0A F5 04 
B7 47 00 00 93 87 47 ED 03 A7 07 00 83 A6 89 00 
B3 84 84 40 93 E4 14 00 33 04 87 40 13 05 09 00 
23 A2 96 00 23 A0 87 00 EF F0 8F 9A 83 20 C1 01 
03 24 81 01 83 24 41 01 03 29 01 01 83 29 C1 00 
03 2A 81 00 13 05 10 00 13 01 01 02 67 80 00 00 
93 05 00 00 13 05 09 00 EF F0 4F EF 03 A7 89 00 
93 06 F0 00 B3 07 E5 40 E3 DC F6 F4 B7 46 00 00 
83 A6 06 EA 93 E7 17 00 23 22 F7 00 33 05 D5 40 
B7 46 00 00 23 AA A6 EC 6F F0 9F F3 63 8A 05 12 
13 01 01 FF 23 24 81 00 23 22 91 00 13 84 05 00 
93 04 05 00 23 26 11 00 EF F0 4F 92 03 28 C4 FF 
13 07 84 FF B7 45 00 00 93 77 E8 FF 33 06 F7 00 
93 85 05 A9 83 26 46 00 03 A5 85 00 93 F6 C6 FF 
63 0A C5 1A 23 22 D6 00 13 78 18 00 33 05 D6 00 
63 10 08 0A 03 23 84 FF 03 28 45 00 37 45 00 00 
33 07 67 40 83 28 87 00 13 05 85 A9 B3 87 67 00 
13 78 18 00 63 80 A8 14 03 23 C7 00 23 A6 68 00 
23 24 13 01 63 04 08 1E 93 E6 17 00 23 22 D7 00 
23 20 F6 00 93 06 F0 1F 63 E8 F6 0A 93 F6 87 FF 
93 86 86 00 03 A5 45 00 B3 86 D5 00 03 A6 06 00 
13 D8 57 00 93 07 10 00 B3 97 07 01 B3 E7 A7 00 
13 85 86 FF 23 26 A7 00 23 24 C7 00 23 A2 F5 00 
23 A0 E6 00 23 26 E6 00 03 24 81 00 83 20 C1 00 
13 85 04 00 83 24 41 00 13 01 01 01 6F F0 4F 85 
03 25 45 00 13 75 15 00 63 1E 05 02 37 45 00 00 
B3 87 D7 00 13 05 85 A9 83 26 86 00 93 E8 17 00 
33 08 F7 00 63 88 A6 16 03 26 C6 00 23 A6 C6 00 
23 24 D6 00 23 22 17 01 23 20 F8 00 6F F0 9F F6 
67 80 00 00 93 E6 17 00 23 2E D4 FE 23 20 F6 00 
93 06 F0 1F E3 FC F6 F4 93 D6 97 00 13 06 40 00 
63 6C D6 0E 93 D6 67 00 13 88 96 03 13 86 86 03 
13 18 38 00 33 88 05 01 83 26 08 00 13 08 88 FF 
63 08 D8 12 03 A6 46 00 13 76 C6 FF 63 F6 C7 00 
83 A6 86 00 E3 18 D8 FE 03 A8 C6 00 23 26 07 01 
23 24 D7 00 03 24 81 00 83 20 C1 00 23 24 E8 00 
13 85 04 00 83 24 41 00 23 A6 E6 00 13 01 01 01 
6F E0 1F F9 63 16 08 14 83 25 C6 00 03 26 86 00 
B3 87 F6 00 03 24 81 00 23 26 B6 00 23 A4 C5 00 
93 E6 17 00 83 20 C1 00 23 22 D7 00 13 85 04 00 
33 07 F7 00 83 24 41 00 23 20 F7 00 13 01 01 01 
6F E0 1F F5 13 78 18 00 B3 87 D7 00 63 10 08 02 
03 25 84 FF 33 07 A7 40 83 26 C7 00 03 26 87 00 
B3 87 A7 00 23 26 D6 00 23 A4 C6 00 B7 46 00 00 
13 E6 17 00 83 A6 46 EA 23 22 C7 00 23 A4 E5 00 
E3 E4 D7 EA B7 47 00 00 83 A5 87 F0 13 85 04 00 
EF F0 DF C7 6F F0 5F E9 13 06 40 01 63 74 D6 02 
13 06 40 05 63 64 D6 06 93 D6 C7 00 13 88 F6 06 
13 86 E6 06 13 18 38 00 6F F0 DF EF B3 87 D7 00 
6F F0 9F E9 13 88 C6 05 13 86 B6 05 13 18 38 00 
6F F0 5F EE 23 AA E5 00 23 A8 E5 00 23 26 A7 00 
23 24 A7 00 23 22 17 01 23 20 F8 00 6F F0 DF E3 
03 A5 45 00 13 56 26 40 93 07 10 00 33 96 C7 00 
33 66 A6 00 23 A2 C5 00 6F F0 5F ED 13 06 40 15 
63 6C D6 00 93 D6 F7 00 13 88 86 07 13 86 76 07 
13 18 38 00 6F F0 1F E9 13 06 40 55 63 6C D6 00 
93 D6 27 01 13 88 D6 07 13 86 C6 07 13 18 38 00 
6F F0 5F E7 13 08 80 3F 13 06 E0 07 6F F0 9F E6 
93 E6 17 00 23 22 D7 00 23 20 F6 00 6F F0 DF DC 
13 01 01 FF 13 87 05 00 23 24 81 00 23 22 91 00 
93 05 06 00 13 04 05 00 B7 44 00 00 13 86 06 00 
13 05 07 00 23 26 11 00 23 AE 04 EE EF 00 40 69 
93 07 F0 FF 63 0C F5 00 83 20 C1 00 03 24 81 00 
83 24 41 00 13 01 01 01 67 80 00 00 83 A7 C4 EF 
E3 84 07 FE 83 20 C1 00 23 20 F4 00 03 24 81 00 
83 24 41 00 13 01 01 01 67 80 00 00 13 01 01 F9 
23 24 81 06 13 84 05 00 83 95 E5 00 23 22 91 06 
23 20 21 07 23 26 11 06 93 04 06 00 13 89 06 00 
63 CA 05 04 13 06 81 00 EF 00 40 41 63 44 05 04 
03 27 C1 00 B7 F7 00 00 83 20 C1 06 B3 F7 E7 00 
37 E7 FF FF B3 87 E7 00 03 24 81 06 93 B7 17 00 
23 20 F9 00 93 07 00 40 23 A0 F4 00 37 15 00 00 
83 24 41 06 03 29 01 06 13 05 05 80 13 01 01 07 
67 80 00 00 83 57 C4 00 23 20 09 00 93 F7 07 08 
63 84 07 02 83 20 C1 06 03 24 81 06 93 07 00 04 
23 A0 F4 00 03 29 01 06 83 24 41 06 13 05 00 00 
13 01 01 07 67 80 00 00 83 20 C1 06 03 24 81 06 
93 07 00 40 23 A0 F4 00 03 29 01 06 83 24 41 06 
13 05 00 00 13 01 01 07 67 80 00 00 83 D7 C5 00 
13 01 01 FE 23 2C 81 00 23 2E 11 00 23 2A 91 00 
23 28 21 01 93 F7 27 00 13 84 05 00 63 88 07 02 
93 87 35 04 23 A0 F5 00 23 A8 F5 00 93 07 10 00 
23 AA F5 00 83 20 C1 01 03 24 81 01 83 24 41 01 
03 29 01 01 13 01 01 02 67 80 00 00 93 06 C1 00 
13 06 81 00 93 04 05 00 EF F0 5F ED 83 25 81 00 
13 09 05 00 13 85 04 00 EF E0 8F AD 83 17 C4 00 
63 06 05 04 13 07 C0 69 23 AE E4 02 03 27 81 00 
83 26 C1 00 93 E7 07 08 23 16 F4 00 23 20 A4 00 
23 28 A4 00 23 2A E4 00 63 98 06 04 B3 E7 27 01 
83 20 C1 01 23 16 F4 00 03 24 81 01 83 24 41 01 
03 29 01 01 13 01 01 02 67 80 00 00 13 F7 07 20 
E3 1A 07 F6 93 F7 C7 FF 93 E7 27 00 13 07 34 04 
23 16 F4 00 93 07 10 00 23 20 E4 00 23 28 E4 00 
23 2A F4 00 6F F0 1F F5 83 15 E4 00 13 85 04 00 
EF 00 40 2E 63 16 05 00 83 17 C4 00 6F F0 1F FA 
03 57 C4 00 13 77 C7 FF 13 67 17 00 93 17 07 01 
93 D7 07 41 6F F0 9F F8 13 01 01 FF 13 87 05 00 
23 24 81 00 23 22 91 00 93 05 06 00 13 04 05 00 
B7 44 00 00 13 86 06 00 13 05 07 00 23 26 11 00 
23 AE 04 EE EF 00 C0 48 93 07 F0 FF 63 0C F5 00 
83 20 C1 00 03 24 81 00 83 24 41 00 13 01 01 01 
67 80 00 00 83 A7 C4 EF E3 84 07 FE 83 20 C1 00 
23 20 F4 00 03 24 81 00 83 24 41 00 13 01 01 01 
67 80 00 00 13 01 01 FF 23 24 81 00 13 84 05 00 
83 A5 05 00 23 22 91 00 23 26 11 00 93 04 05 00 
63 84 05 00 EF F0 1F FE 93 05 04 00 03 24 81 00 
83 20 C1 00 13 85 04 00 83 24 41 00 13 01 01 01 
6F F0 DF 9E B7 47 00 00 83 A7 C7 E9 63 80 A7 10 
83 25 C5 04 13 01 01 FE 23 2A 91 00 23 2E 11 00 
23 2C 81 00 23 28 21 01 23 26 31 01 93 04 05 00 
63 80 05 04 13 09 00 00 93 09 00 08 B3 87 25 01 
03 A4 07 00 63 0E 04 00 93 05 04 00 03 24 04 00 
13 85 04 00 EF F0 9F 99 E3 18 04 FE 83 A5 C4 04 
13 09 49 00 E3 1C 39 FD 13 85 04 00 EF F0 1F 98 
83 A5 04 04 63 86 05 00 13 85 04 00 EF F0 1F 97 
03 A4 84 14 63 00 04 02 13 89 C4 14 63 0C 24 01 
93 05 04 00 03 24 04 00 13 85 04 00 EF F0 1F 95 
E3 18 89 FE 83 A5 44 05 63 86 05 00 13 85 04 00 
EF F0 DF 93 83 A7 84 03 63 8C 07 02 83 A7 C4 03 
13 85 04 00 E7 80 07 00 83 A5 04 2E 63 82 05 02 
03 24 81 01 83 20 C1 01 03 29 01 01 83 29 C1 00 
13 85 04 00 83 24 41 01 13 01 01 02 6F F0 9F ED 
83 20 C1 01 03 24 81 01 83 24 41 01 03 29 01 01 
83 29 C1 00 13 01 01 02 67 80 00 00 67 80 00 00 
B7 37 00 00 03 A7 07 66 83 27 87 14 63 8C 07 04 
03 A7 47 00 13 08 F0 01 63 4E E8 06 13 18 27 00 
63 06 05 02 33 83 07 01 23 24 C3 08 83 A8 87 18 
13 06 10 00 33 16 E6 00 B3 E8 C8 00 23 A4 17 19 
23 24 D3 10 93 06 20 00 63 04 D5 02 13 07 17 00 
23 A2 E7 00 B3 87 07 01 23 A4 B7 00 13 05 00 00 
67 80 00 00 93 07 C7 14 23 24 F7 14 6F F0 5F FA 
83 A6 C7 18 13 07 17 00 23 A2 E7 00 33 E6 C6 00 
23 A6 C7 18 B3 87 07 01 23 A4 B7 00 13 05 00 00 
67 80 00 00 13 05 F0 FF 67 80 00 00 13 01 01 FF 
13 87 05 00 23 24 81 00 23 22 91 00 13 04 05 00 
B7 44 00 00 93 05 06 00 13 05 07 00 23 26 11 00 
23 AE 04 EE EF 00 C0 13 93 07 F0 FF 63 0C F5 00 
83 20 C1 00 03 24 81 00 83 24 41 00 13 01 01 01 
67 80 00 00 83 A7 C4 EF E3 84 07 FE 83 20 C1 00 
23 20 F4 00 03 24 81 00 83 24 41 00 13 01 01 01 
67 80 00 00 13 01 01 FF 23 24 81 00 23 22 91 00 
13 04 05 00 B7 44 00 00 13 85 05 00 23 26 11 00 
23 AE 04 EE EF 00 C0 14 93 07 F0 FF 63 0C F5 00 
83 20 C1 00 03 24 81 00 83 24 41 00 13 01 01 01 
67 80 00 00 83 A7 C4 EF E3 84 07 FE 83 20 C1 00 
23 20 F4 00 03 24 81 00 83 24 41 00 13 01 01 01 
67 80 00 00 13 01 01 FF 23 26 11 00 23 24 81 00 
93 05 00 00 13 06 00 00 93 06 00 00 13 07 00 00 
93 07 00 00 93 08 90 03 73 00 00 00 13 04 05 00 
63 4C 05 00 83 20 C1 00 13 05 04 00 03 24 81 00 
13 01 01 01 67 80 00 00 33 04 80 40 EF 00 80 2E 
23 20 85 00 13 04 F0 FF 6F F0 DF FD 93 05 00 00 
13 06 00 00 93 06 00 00 13 07 00 00 93 07 00 00 
93 08 D0 05 73 00 00 00 63 44 05 00 6F 00 00 00 
13 01 01 FF 23 24 81 00 13 04 05 00 23 26 11 00 
33 04 80 40 EF 00 00 2A 23 20 85 00 6F 00 00 00 
13 01 01 F7 23 22 91 08 23 26 11 08 93 84 05 00 
23 24 81 08 93 05 01 00 13 06 00 00 93 06 00 00 
13 07 00 00 93 07 00 00 93 08 00 05 73 00 00 00 
13 04 05 00 63 44 05 02 13 85 04 00 93 05 01 00 
EF 00 00 1B 83 20 C1 08 13 05 04 00 03 24 81 08 
83 24 41 08 13 01 01 09 67 80 00 00 33 04 80 40 
EF 00 40 23 23 20 85 00 13 04 F0 FF 6F F0 DF FC 
13 01 01 F9 93 05 81 00 23 26 11 06 EF F0 5F F8 
93 07 F0 FF 63 0E F5 00 03 25 C1 00 83 20 C1 06 
13 55 D5 00 13 75 15 00 13 01 01 07 67 80 00 00 
83 20 C1 06 13 05 00 00 13 01 01 07 67 80 00 00 
13 01 01 FF 23 26 11 00 23 24 81 00 93 06 00 00 
13 07 00 00 93 07 00 00 93 08 E0 03 73 00 00 00 
13 04 05 00 63 4C 05 00 83 20 C1 00 13 05 04 00 
03 24 81 00 13 01 01 01 67 80 00 00 33 04 80 40 
EF 00 40 1A 23 20 85 00 13 04 F0 FF 6F F0 DF FD 
13 01 01 FF 23 26 11 00 23 24 81 00 93 06 00 00 
13 07 00 00 93 07 00 00 93 08 F0 03 73 00 00 00 
13 04 05 00 63 4C 05 00 83 20 C1 00 13 05 04 00 
03 24 81 00 13 01 01 01 67 80 00 00 33 04 80 40 
EF 00 40 15 23 20 85 00 13 04 F0 FF 6F F0 DF FD 
37 43 00 00 83 27 C3 F0 13 01 01 FF 23 26 11 00 
13 08 05 00 63 98 07 02 13 05 00 00 93 05 00 00 
13 06 00 00 93 06 00 00 13 07 00 00 93 08 60 0D 
73 00 00 00 13 07 F0 FF 93 07 05 00 63 04 E5 04 
23 26 A3 F0 33 05 F8 00 93 05 00 00 13 06 00 00 
93 06 00 00 13 07 00 00 93 07 00 00 93 08 60 0D 
73 00 00 00 83 27 C3 F0 33 08 F8 00 63 1C 05 01 
83 20 C1 00 23 26 A3 F0 13 85 07 00 13 01 01 01 
67 80 00 00 EF 00 00 0C 83 20 C1 00 93 07 C0 00 
23 20 F5 00 13 05 F0 FF 13 01 01 01 67 80 00 00 
13 01 01 FF 83 A3 45 01 83 A2 85 01 83 AF C5 01 
03 AF 05 02 83 AE 05 03 03 AE 05 04 03 A3 85 03 
03 A8 85 04 83 A8 C5 04 03 A6 85 05 23 26 81 00 
23 24 91 00 03 A4 05 01 83 A4 85 00 23 22 21 01 
03 A9 05 00 83 A6 C5 05 03 A7 85 06 83 A7 C5 06 
23 10 25 01 23 11 95 00 23 22 85 00 23 14 75 00 
23 15 55 00 23 16 F5 01 23 17 E5 01 23 28 D5 01 
23 24 C5 05 23 22 65 04 23 2C 05 01 23 2E 15 01 
23 24 C5 02 23 26 D5 02 03 24 C1 00 23 2C E5 02 
23 2E F5 02 83 24 81 00 03 29 41 00 13 01 01 01 
67 80 00 00 B7 47 00 00 03 A5 C7 E9 67 80 00 00 
13 01 01 FC 23 2C 81 02 23 2A 91 02 23 28 21 03 
23 26 31 03 23 24 41 03 23 2E 11 02 B7 07 00 02 
13 07 00 05 37 35 00 00 23 80 E7 00 13 05 45 60 
EF D0 4F 82 13 04 F0 FF 37 3A 00 00 37 39 00 00 
B7 34 00 00 93 09 A0 00 13 06 10 01 93 05 8A 64 
13 05 C1 00 EF C0 9F D3 93 57 84 01 93 06 01 02 
93 F7 F7 00 B3 87 F6 00 83 C7 C7 FE 13 57 C4 01 
33 87 E6 00 03 47 C7 FE A3 02 F1 00 93 57 04 01 
93 F7 F7 0F 23 02 E1 00 13 D7 47 00 93 F7 F7 00 
B3 87 F6 00 83 C7 C7 FE 33 87 E6 00 03 47 C7 FE 
A3 03 F1 00 93 57 84 00 93 F7 F7 0F 23 03 E1 00 
13 D7 47 00 93 F7 F7 00 B3 87 F6 00 33 87 E6 00 
83 C7 C7 FE 03 47 C7 FE 13 06 20 00 A3 04 F1 00 
93 77 F4 0F 23 04 E1 00 13 D7 47 00 93 F7 F7 00 
33 87 E6 00 B3 87 F6 00 03 47 C7 FE 83 C7 C7 FE 
93 05 49 62 37 05 00 01 23 05 E1 00 A3 05 F1 00 
EF C0 1F B6 13 06 80 00 93 05 41 00 37 05 00 01 
EF C0 1F B5 13 06 20 00 93 85 84 62 37 05 00 01 
13 04 14 00 EF C0 DF B3 E3 10 34 F3 37 35 00 00 
13 05 C5 62 EF C0 1F F2 B7 04 00 01 37 04 00 02 
83 A7 04 00 23 26 F1 00 13 97 07 01 E3 5A 07 FE 
13 06 10 00 93 05 C1 00 37 05 00 01 EF C0 5F B0 
83 47 C1 00 23 00 F4 00 6F F0 9F FD B7 07 00 00 
93 87 07 00 63 86 07 00 13 85 41 1F 6F E0 9F D0 
67 80 00 00 
@00003604
4E 6F 77 20 72 75 6E 6E 69 6E 67 3A 20 43 6F 75 
6E 74 20 66 72 6F 6D 20 2D 31 20 74 6F 20 39 00 
30 78 00 00 0D 0A 00 00 4E 6F 77 20 72 75 6E 6E 
69 6E 67 3A 20 55 41 52 54 20 4C 6F 6F 70 62 61 
63 6B 00 00 30 31 32 33 34 35 36 37 38 39 61 62 
63 64 65 66 00 00 00 00 0A 00 00 00 
@00003660
68 36 00 00 
@00003668
00 00 00 00 54 39 00 00 BC 39 00 00 24 3A 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 01 00 00 00 00 00 00 00 
0E 33 CD AB 34 12 6D E6 EC DE 05 00 0B 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 
90 3A 00 00 90 3A 00 00 98 3A 00 00 98 3A 00 00 
A0 3A 00 00 A0 3A 00 00 A8 3A 00 00 A8 3A 00 00 
B0 3A 00 00 B0 3A 00 00 B8 3A 00 00 B8 3A 00 00 
C0 3A 00 00 C0 3A 00 00 C8 3A 00 00 C8 3A 00 00 
D0 3A 00 00 D0 3A 00 00 D8 3A 00 00 D8 3A 00 00 
E0 3A 00 00 E0 3A 00 00 E8 3A 00 00 E8 3A 00 00 
F0 3A 00 00 F0 3A 00 00 F8 3A 00 00 F8 3A 00 00 
00 3B 00 00 00 3B 00 00 08 3B 00 00 08 3B 00 00 
10 3B 00 00 10 3B 00 00 18 3B 00 00 18 3B 00 00 
20 3B 00 00 20 3B 00 00 28 3B 00 00 28 3B 00 00 
30 3B 00 00 30 3B 00 00 38 3B 00 00 38 3B 00 00 
40 3B 00 00 40 3B 00 00 48 3B 00 00 48 3B 00 00 
50 3B 00 00 50 3B 00 00 58 3B 00 00 58 3B 00 00 
60 3B 00 00 60 3B 00 00 68 3B 00 00 68 3B 00 00 
70 3B 00 00 70 3B 00 00 78 3B 00 00 78 3B 00 00 
80 3B 00 00 80 3B 00 00 88 3B 00 00 88 3B 00 00 
90 3B 00 00 90 3B 00 00 98 3B 00 00 98 3B 00 00 
A0 3B 00 00 A0 3B 00 00 A8 3B 00 00 A8 3B 00 00 
B0 3B 00 00 B0 3B 00 00 B8 3B 00 00 B8 3B 00 00 
C0 3B 00 00 C0 3B 00 00 C8 3B 00 00 C8 3B 00 00 
D0 3B 00 00 D0 3B 00 00 D8 3B 00 00 D8 3B 00 00 
E0 3B 00 00 E0 3B 00 00 E8 3B 00 00 E8 3B 00 00 
F0 3B 00 00 F0 3B 00 00 F8 3B 00 00 F8 3B 00 00 
00 3C 00 00 00 3C 00 00 08 3C 00 00 08 3C 00 00 
10 3C 00 00 10 3C 00 00 18 3C 00 00 18 3C 00 00 
20 3C 00 00 20 3C 00 00 28 3C 00 00 28 3C 00 00 
30 3C 00 00 30 3C 00 00 38 3C 00 00 38 3C 00 00 
40 3C 00 00 40 3C 00 00 48 3C 00 00 48 3C 00 00 
50 3C 00 00 50 3C 00 00 58 3C 00 00 58 3C 00 00 
60 3C 00 00 60 3C 00 00 68 3C 00 00 68 3C 00 00 
70 3C 00 00 70 3C 00 00 78 3C 00 00 78 3C 00 00 
80 3C 00 00 80 3C 00 00 88 3C 00 00 88 3C 00 00 
90 3C 00 00 90 3C 00 00 98 3C 00 00 98 3C 00 00 
A0 3C 00 00 A0 3C 00 00 A8 3C 00 00 A8 3C 00 00 
B0 3C 00 00 B0 3C 00 00 B8 3C 00 00 B8 3C 00 00 
C0 3C 00 00 C0 3C 00 00 C8 3C 00 00 C8 3C 00 00 
D0 3C 00 00 D0 3C 00 00 D8 3C 00 00 D8 3C 00 00 
E0 3C 00 00 E0 3C 00 00 E8 3C 00 00 E8 3C 00 00 
F0 3C 00 00 F0 3C 00 00 F8 3C 00 00 F8 3C 00 00 
00 3D 00 00 00 3D 00 00 08 3D 00 00 08 3D 00 00 
10 3D 00 00 10 3D 00 00 18 3D 00 00 18 3D 00 00 
20 3D 00 00 20 3D 00 00 28 3D 00 00 28 3D 00 00 
30 3D 00 00 30 3D 00 00 38 3D 00 00 38 3D 00 00 
40 3D 00 00 40 3D 00 00 48 3D 00 00 48 3D 00 00 
50 3D 00 00 50 3D 00 00 58 3D 00 00 58 3D 00 00 
60 3D 00 00 60 3D 00 00 68 3D 00 00 68 3D 00 00 
70 3D 00 00 70 3D 00 00 78 3D 00 00 78 3D 00 00 
80 3D 00 00 80 3D 00 00 88 3D 00 00 88 3D 00 00 
90 3D 00 00 90 3D 00 00 98 3D 00 00 98 3D 00 00 
A0 3D 00 00 A0 3D 00 00 A8 3D 00 00 A8 3D 00 00 
B0 3D 00 00 B0 3D 00 00 B8 3D 00 00 B8 3D 00 00 
C0 3D 00 00 C0 3D 00 00 C8 3D 00 00 C8 3D 00 00 
D0 3D 00 00 D0 3D 00 00 D8 3D 00 00 D8 3D 00 00 
E0 3D 00 00 E0 3D 00 00 E8 3D 00 00 E8 3D 00 00 
F0 3D 00 00 F0 3D 00 00 F8 3D 00 00 F8 3D 00 00 
00 3E 00 00 00 3E 00 00 08 3E 00 00 08 3E 00 00 
10 3E 00 00 10 3E 00 00 18 3E 00 00 18 3E 00 00 
20 3E 00 00 20 3E 00 00 28 3E 00 00 28 3E 00 00 
30 3E 00 00 30 3E 00 00 38 3E 00 00 38 3E 00 00 
40 3E 00 00 40 3E 00 00 48 3E 00 00 48 3E 00 00 
50 3E 00 00 50 3E 00 00 58 3E 00 00 58 3E 00 00 
60 3E 00 00 60 3E 00 00 68 3E 00 00 68 3E 00 00 
70 3E 00 00 70 3E 00 00 78 3E 00 00 78 3E 00 00 
80 3E 00 00 80 3E 00 00 88 3E 00 00 88 3E 00 00 
00 00 00 00 68 36 00 00 FF FF FF FF 00 00 02 00 
@00003EA8
00 00 00 00 
@00003EAC
64 00 00 00 
@00003EB0
B8 00 00 00 
@00003EB4
EC 35 00 00 
