@00000000
17 11 00 00 13 01 01 00 6F 00 00 02 63 5C C0 00 
33 86 C5 00 83 C7 05 00 93 85 15 00 23 00 F5 00 
E3 9A C5 FE 67 80 00 00 13 01 01 FF 23 26 11 00 
EF 00 40 00 B7 07 00 02 13 07 50 05 23 80 E7 00 
B7 07 00 01 13 07 80 04 23 80 E7 00 13 07 50 06 
23 80 E7 00 13 07 C0 06 23 80 E7 00 23 80 E7 00 
93 06 F0 06 23 80 D7 00 13 06 C0 02 23 80 C7 00 
13 06 00 02 23 80 C7 00 13 06 70 05 23 80 C7 00 
23 80 D7 00 93 06 20 07 23 80 D7 00 23 80 E7 00 
13 07 40 06 23 80 E7 00 13 07 10 02 23 80 E7 00 
13 07 D0 00 23 80 E7 00 13 07 A0 00 23 80 E7 00 
23 80 07 00 6F 00 00 00 
