@00000000
17 11 00 00 13 01 01 00 6F 00 40 00 13 01 01 FF 
23 26 11 00 EF 00 40 00 93 05 80 04 13 06 80 05 
37 07 00 01 93 86 05 00 83 27 47 00 93 D7 07 01 
E3 8C 07 FE 83 C7 06 00 93 86 16 00 23 00 F7 00 
E3 94 C6 FE 6F F0 1F FE 
@00000048
48 65 6C 6C 6F 2C 20 57 6F 72 6C 64 21 0D 0A 00 
