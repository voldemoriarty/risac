@00000000
17 11 00 00 13 01 01 00 6F 00 C0 02 63 52 C0 02 
33 87 C5 00 83 27 45 00 93 D7 07 01 E3 8C 07 FE 
83 C7 05 00 93 85 15 00 23 00 F5 00 E3 94 E5 FE 
67 80 00 00 13 01 01 FF 23 26 11 00 EF 00 40 00 
93 07 00 0E 03 A6 07 02 83 A6 47 02 03 A7 87 02 
03 AF 07 00 83 AE 47 00 03 AE 87 00 03 A3 C7 00 
83 A8 07 01 03 A8 47 01 03 A5 87 01 83 A5 C7 01 
83 C7 C7 02 B7 0F 00 02 93 02 00 05 13 01 01 FD 
23 80 5F 00 23 20 C1 02 23 22 D1 02 23 24 E1 02 
23 20 E1 01 23 22 D1 01 23 24 C1 01 23 26 61 00 
23 28 11 01 23 2A 01 01 23 2C A1 00 23 2E B1 00 
23 06 F1 02 93 06 01 00 13 06 D1 02 37 07 00 01 
83 27 47 00 93 D7 07 01 E3 8C 07 FE 83 C7 06 00 
93 86 16 00 23 00 F7 00 E3 94 C6 FE 6F 00 00 00 
@000000E0
48 6F 77 64 79 20 66 72 69 65 6E 64 2C 20 68 6F 
77 20 67 6F 65 73 20 74 68 65 20 68 75 6E 74 20 
66 6F 72 20 73 6F 75 6C 73 3F 0D 0A 00 00 00 00 
