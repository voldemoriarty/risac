@00000000
17 11 00 00 13 01 01 00 6F 00 00 03 93 07 00 00 
B7 06 00 01 03 A7 46 00 13 57 07 01 E3 0C 07 FE 
33 07 F5 00 03 47 07 00 93 87 17 00 23 80 E6 00 
E3 92 B7 FE 67 80 00 00 13 01 01 FC 23 2C 81 02 
23 2A 91 02 23 28 21 03 23 26 31 03 23 24 41 03 
23 2E 11 02 B7 07 00 02 13 07 00 05 23 80 E7 00 
93 05 20 02 13 05 C0 1A EF F0 5F FA 13 04 F0 FF 
93 09 A0 00 13 06 10 01 93 05 80 1F 13 05 C1 00 
EF 00 80 10 93 57 84 01 93 06 01 02 93 F7 F7 00 
B3 87 F6 00 83 C7 C7 FE 13 57 C4 01 33 87 E6 00 
03 47 C7 FE A3 02 F1 00 93 57 04 01 93 F7 F7 0F 
23 02 E1 00 13 D7 47 00 93 F7 F7 00 B3 87 F6 00 
83 C7 C7 FE 33 87 E6 00 03 47 C7 FE A3 03 F1 00 
93 57 84 00 93 F7 F7 0F 23 03 E1 00 13 D7 47 00 
93 F7 F7 00 B3 87 F6 00 33 87 E6 00 83 C7 C7 FE 
03 47 C7 FE 93 05 20 00 A3 04 F1 00 93 77 F4 0F 
23 04 E1 00 13 D7 47 00 93 F7 F7 00 33 87 E6 00 
B3 87 F6 00 03 47 C7 FE 83 C7 C7 FE 13 05 00 1D 
23 05 E1 00 A3 05 F1 00 EF F0 5F EE 93 05 80 00 
13 05 41 00 EF F0 9F ED 93 05 20 00 13 05 40 1D 
13 04 14 00 EF F0 9F EC E3 16 34 F3 93 05 D0 01 
13 05 80 1D EF F0 9F EB B7 04 00 01 37 04 00 02 
83 A7 04 00 23 26 F1 00 13 97 07 01 E3 5A 07 FE 
93 05 10 00 13 05 C1 00 EF F0 5F E9 83 47 C1 00 
23 00 F4 00 6F F0 DF FD 93 07 00 00 63 94 C7 00 
67 80 00 00 33 87 F5 00 83 46 07 00 33 07 F5 00 
93 87 17 00 23 00 D7 00 6F F0 5F FE 
@000001AC
4E 6F 77 20 72 75 6E 6E 69 6E 67 3A 20 43 6F 75 
6E 74 20 66 72 6F 6D 20 2D 31 20 74 6F 20 39 0D 
0A 00 00 00 30 78 00 00 0D 0A 00 00 4E 6F 77 20 
72 75 6E 6E 69 6E 67 3A 20 55 41 52 54 20 4C 6F 
6F 70 62 61 63 6B 0D 0A 00 00 00 00 30 31 32 33 
34 35 36 37 38 39 61 62 63 64 65 66 00 00 00 00 
