@00000000
17 11 00 00 13 01 01 00 6F 00 00 10 63 52 C0 02 
33 87 C5 00 83 27 45 00 93 D7 07 01 E3 8C 07 FE 
83 C7 05 00 93 85 15 00 23 00 F5 00 E3 94 E5 FE 
67 80 00 00 93 07 80 28 03 CE 07 01 03 AF 87 00 
83 AE C7 00 83 A2 07 00 83 AF 47 00 13 D7 05 01 
93 D7 85 00 13 01 01 FE 93 F6 F5 0F 13 77 F7 0F 
93 F7 F7 0F 13 D6 85 01 23 0E C1 01 13 53 47 00 
13 0E 01 02 93 D8 47 00 13 D8 46 00 93 D5 C5 01 
13 76 F6 00 13 77 F7 00 93 F7 F7 00 93 F6 F6 00 
23 26 51 00 23 28 F1 01 23 2A E1 01 23 2C D1 01 
B3 05 BE 00 33 06 CE 00 33 07 EE 00 B3 07 FE 00 
33 03 6E 00 B3 08 1E 01 33 08 0E 01 B3 06 DE 00 
03 CF C5 FE 83 4E C6 FE 03 4E C3 FE 03 C6 C7 FE 
03 43 C7 FE 83 C5 C8 FE 03 47 C8 FE 83 C7 C6 FE 
23 00 E5 01 A3 00 D5 01 23 01 C5 01 A3 01 65 00 
23 02 B5 00 A3 02 C5 00 23 03 E5 00 A3 03 F5 00 
13 01 01 02 67 80 00 00 13 01 01 FF 23 26 11 00 
EF 00 40 00 13 01 01 FC 93 07 80 28 23 2E 11 02 
37 07 00 02 83 A0 07 00 83 A3 47 00 83 A2 87 00 
83 AF C7 00 03 CF 07 01 23 2C 81 02 23 2A 91 02 
23 28 21 03 23 26 31 03 23 24 41 03 23 22 51 03 
93 06 00 05 B7 17 00 00 23 00 D7 00 93 87 D7 A0 
37 07 00 01 B7 05 FF FF 37 06 01 FF 23 14 F1 00 
13 05 F0 0F 93 0E A1 00 93 85 F5 0F 13 06 F6 FF 
13 08 F7 FF 13 0E 00 03 13 03 80 07 93 08 00 10 
23 26 11 00 93 07 01 02 93 56 85 00 23 28 71 00 
23 2A 51 00 23 2C F1 01 23 0E E1 01 B3 86 D7 00 
13 74 F5 0F 83 47 C1 00 83 CA C6 FE 93 54 44 00 
13 09 01 02 B3 04 99 00 93 86 07 00 13 89 07 00 
83 C9 C4 FE B3 F7 B7 00 93 04 01 02 13 74 F4 00 
33 84 84 00 13 9A 86 00 93 9A 8A 00 93 86 07 00 
83 44 C4 FE B3 E7 57 01 B3 E6 46 01 13 04 09 00 
93 99 09 01 B3 F7 C7 00 13 19 09 01 B3 F6 C6 00 
B3 E7 37 01 B3 E6 26 01 93 94 84 01 B3 F7 07 01 
13 14 84 01 B3 F6 06 01 B3 E7 97 00 B3 E6 86 00 
23 20 D1 00 23 22 F1 00 83 27 47 00 93 D7 07 01 
E3 8C 07 FE 23 00 C7 01 83 27 47 00 93 D7 07 01 
E3 8C 07 FE 23 00 67 00 93 06 01 00 83 27 47 00 
93 D7 07 01 E3 8C 07 FE 83 C7 06 00 93 86 16 00 
23 00 F7 00 E3 94 DE FE 63 06 15 01 13 05 00 10 
6F F0 1F F1 6F 00 00 00 
@00000288
30 31 32 33 34 35 36 37 38 39 61 62 63 64 65 66 
00 00 00 00 
