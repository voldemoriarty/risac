@00000000
17 11 00 00 13 01 01 00 6F 00 40 00 13 01 01 FF 
23 26 11 00 EF 00 40 00 93 07 80 08 03 A6 87 00 
83 A6 C7 00 03 A7 07 01 03 A5 07 00 83 A5 47 00 
83 D7 47 01 37 08 00 02 93 08 50 05 13 01 01 FE 
23 00 18 01 23 28 C1 00 23 2A D1 00 23 2C E1 00 
23 24 A1 00 23 26 B1 00 23 1E F1 00 93 06 81 00 
13 06 E1 01 37 07 00 01 83 27 47 00 93 D7 07 01 
E3 8C 07 FE 83 C7 06 00 93 86 16 00 23 00 F7 00 
E3 94 C6 FE 6F 00 00 00 
@00000088
48 6F 77 64 79 20 64 6F 77 64 79 20 64 6F 6F 20 
64 61 61 0D 0A 00 00 00 
