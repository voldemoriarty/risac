@00000000
17 11 00 00 13 01 01 00 6F 00 80 27 63 52 C0 02 
33 87 C5 00 83 27 45 00 93 D7 07 01 E3 8C 07 FE 
83 C7 05 00 93 85 15 00 23 00 F5 00 E3 94 E5 FE 
67 80 00 00 93 07 40 42 03 CE 07 01 03 AF 87 00 
83 AE C7 00 83 A2 07 00 83 AF 47 00 13 D7 05 01 
93 D7 85 00 13 01 01 FE 93 F6 F5 0F 13 77 F7 0F 
93 F7 F7 0F 13 D6 85 01 23 0E C1 01 13 53 47 00 
13 0E 01 02 93 D8 47 00 13 D8 46 00 93 D5 C5 01 
13 76 F6 00 13 77 F7 00 93 F7 F7 00 93 F6 F6 00 
23 26 51 00 23 28 F1 01 23 2A E1 01 23 2C D1 01 
B3 05 BE 00 33 06 CE 00 33 07 EE 00 B3 07 FE 00 
33 03 6E 00 B3 08 1E 01 33 08 0E 01 B3 06 DE 00 
03 CF C5 FE 83 4E C6 FE 03 4E C3 FE 03 C6 C7 FE 
03 43 C7 FE 83 C5 C8 FE 03 47 C8 FE 83 C7 C6 FE 
23 00 E5 01 A3 00 D5 01 23 01 C5 01 A3 01 65 00 
23 02 B5 00 A3 02 C5 00 23 03 E5 00 A3 03 F5 00 
13 01 01 02 67 80 00 00 93 07 40 42 83 C6 07 01 
83 AE 47 00 03 AE 87 00 03 A3 C7 00 03 AF 07 00 
93 D7 85 00 13 01 01 FE 93 F7 F7 0F 23 0E D1 00 
13 D6 85 01 93 D8 47 00 93 06 01 02 93 F7 F7 00 
B3 88 16 01 13 D7 05 01 B3 86 F6 00 13 D8 C5 01 
93 07 01 02 13 76 F6 00 23 26 E1 01 23 28 D1 01 
23 2A C1 01 23 2C 61 00 13 77 F7 0F 33 88 07 01 
33 86 C7 00 93 F5 F5 0F 83 C7 C8 FE 83 CE C6 FE 
03 4E C6 FE 83 46 C8 FE 93 D8 45 00 13 08 01 02 
13 56 47 00 B3 08 18 01 33 06 C8 00 37 08 FF FF 
13 08 F8 0F 03 C3 C8 FE 93 F5 F5 00 83 48 C6 FE 
13 76 F7 00 33 F7 07 01 93 07 01 02 B3 87 B7 00 
93 05 01 02 B3 F6 06 01 33 86 C5 00 93 9E 8E 00 
13 1E 8E 00 B7 05 01 FF 93 85 F5 FF 03 C8 C7 FE 
03 46 C6 FE B3 67 D7 01 33 E7 C6 01 B3 F7 B7 00 
33 77 B7 00 13 13 03 01 93 98 08 01 B7 06 00 01 
93 86 F6 FF B3 E7 67 00 33 67 17 01 93 15 88 01 
B3 F7 D7 00 13 16 86 01 33 77 D7 00 B3 E7 B7 00 
33 67 C7 00 23 22 E1 00 23 24 F1 00 83 27 45 00 
93 D7 07 01 E3 8C 07 FE 93 07 00 03 23 00 F5 00 
83 27 45 00 93 D7 07 01 E3 8C 07 FE 93 07 80 07 
23 00 F5 00 13 07 41 00 93 06 C1 00 83 27 45 00 
93 D7 07 01 E3 8C 07 FE 83 47 07 00 13 07 17 00 
23 00 F5 00 E3 94 E6 FE 13 01 01 02 67 80 00 00 
13 01 01 FF 23 26 11 00 EF 00 40 00 13 01 01 FB 
93 07 40 42 23 26 11 04 23 24 81 04 23 22 91 04 
03 A4 47 00 83 A4 07 00 83 A0 87 00 83 A3 C7 00 
83 C2 07 01 23 20 21 05 23 2E 31 03 23 2C 41 03 
23 2A 51 03 23 28 61 03 23 26 71 03 37 07 00 01 
B7 07 00 02 93 06 00 05 B7 05 FF FF 37 06 01 FF 
23 80 D7 00 13 05 F0 0F 93 0F C1 00 93 85 F5 0F 
13 06 F6 FF 13 08 F7 FF 13 0F 00 03 93 0E 80 07 
13 0E D0 00 13 03 A0 00 93 08 00 10 23 26 91 00 
93 07 01 02 93 56 85 00 23 28 81 00 23 2A 11 00 
23 2C 71 00 23 0E 51 00 B3 86 D7 00 13 79 F5 0F 
83 47 C1 00 83 CB C6 FE 93 59 49 00 13 0A 01 02 
B3 09 3A 01 93 86 07 00 03 CA C9 FE 93 0A 01 02 
93 89 07 00 13 79 F9 00 B3 F7 B7 00 33 89 2A 01 
13 9B 86 00 93 9B 8B 00 93 86 07 00 83 4A C9 FE 
B3 E7 77 01 B3 E6 66 01 13 89 09 00 13 1A 0A 01 
93 99 09 01 B3 F7 C7 00 B3 F6 C6 00 B3 E6 36 01 
B3 E7 47 01 93 99 8A 01 B3 F7 07 01 13 19 89 01 
B3 F6 06 01 B3 E7 37 01 B3 E6 26 01 23 22 D1 00 
23 24 F1 00 83 27 47 00 93 D7 07 01 E3 8C 07 FE 
23 00 E7 01 83 27 47 00 93 D7 07 01 E3 8C 07 FE 
23 00 D7 01 93 06 41 00 83 27 47 00 93 D7 07 01 
E3 8C 07 FE 83 C7 06 00 93 86 16 00 23 00 F7 00 
E3 94 DF FE 83 27 47 00 93 D7 07 01 E3 8C 07 FE 
23 00 C7 01 83 27 47 00 93 D7 07 01 E3 8C 07 FE 
23 00 67 00 63 06 15 01 13 05 00 10 6F F0 1F EF 
6F 00 00 00 
@00000424
30 31 32 33 34 35 36 37 38 39 61 62 63 64 65 66 
00 00 00 00 
