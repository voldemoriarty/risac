// soc_simple.v

// Generated using ACDS version 19.1 670

`timescale 1 ps / 1 ps
module soc_simple (
		input  wire       clk_clk,       //    clk.clk
		output wire [7:0] leds_export,   //   leds.export
		output wire       locked_export, // locked.export
		input  wire       reset_reset_n  //  reset.reset_n
	);

	wire         pll_50_150_outclk0_clk;                                       // PLL_50_150:outclk_0 -> [jtag_uart:clk, jtag_uart_pipeline_bridge:clk, leds:clk, mm_interconnect_0:PLL_50_150_outclk0_clk, mm_interconnect_1:PLL_50_150_outclk0_clk, mm_interconnect_2:PLL_50_150_outclk0_clk, on_chip_memory:clk, pio_pipeline_bridge:clk, rst_controller:clk, rv32i_core:clk]
	wire  [31:0] rv32i_core_data_master_readdata;                              // mm_interconnect_0:rv32i_core_data_master_readdata -> rv32i_core:avDB_readdata
	wire         rv32i_core_data_master_waitrequest;                           // mm_interconnect_0:rv32i_core_data_master_waitrequest -> rv32i_core:avDB_waitrequest
	wire  [31:0] rv32i_core_data_master_address;                               // rv32i_core:avDB_address -> mm_interconnect_0:rv32i_core_data_master_address
	wire         rv32i_core_data_master_read;                                  // rv32i_core:avDB_read -> mm_interconnect_0:rv32i_core_data_master_read
	wire   [3:0] rv32i_core_data_master_byteenable;                            // rv32i_core:avDB_byteenable -> mm_interconnect_0:rv32i_core_data_master_byteenable
	wire  [31:0] rv32i_core_data_master_writedata;                             // rv32i_core:avDB_writedata -> mm_interconnect_0:rv32i_core_data_master_writedata
	wire         rv32i_core_data_master_write;                                 // rv32i_core:avDB_write -> mm_interconnect_0:rv32i_core_data_master_write
	wire  [31:0] rv32i_core_instruction_master_readdata;                       // mm_interconnect_0:rv32i_core_instruction_master_readdata -> rv32i_core:avIB_readdata
	wire         rv32i_core_instruction_master_waitrequest;                    // mm_interconnect_0:rv32i_core_instruction_master_waitrequest -> rv32i_core:avIB_waitrequest
	wire  [31:0] rv32i_core_instruction_master_address;                        // rv32i_core:avIB_address -> mm_interconnect_0:rv32i_core_instruction_master_address
	wire         rv32i_core_instruction_master_read;                           // rv32i_core:avIB_read -> mm_interconnect_0:rv32i_core_instruction_master_read
	wire  [31:0] mm_interconnect_0_jtag_uart_pipeline_bridge_s0_readdata;      // jtag_uart_pipeline_bridge:s0_readdata -> mm_interconnect_0:jtag_uart_pipeline_bridge_s0_readdata
	wire         mm_interconnect_0_jtag_uart_pipeline_bridge_s0_waitrequest;   // jtag_uart_pipeline_bridge:s0_waitrequest -> mm_interconnect_0:jtag_uart_pipeline_bridge_s0_waitrequest
	wire         mm_interconnect_0_jtag_uart_pipeline_bridge_s0_debugaccess;   // mm_interconnect_0:jtag_uart_pipeline_bridge_s0_debugaccess -> jtag_uart_pipeline_bridge:s0_debugaccess
	wire   [2:0] mm_interconnect_0_jtag_uart_pipeline_bridge_s0_address;       // mm_interconnect_0:jtag_uart_pipeline_bridge_s0_address -> jtag_uart_pipeline_bridge:s0_address
	wire         mm_interconnect_0_jtag_uart_pipeline_bridge_s0_read;          // mm_interconnect_0:jtag_uart_pipeline_bridge_s0_read -> jtag_uart_pipeline_bridge:s0_read
	wire   [3:0] mm_interconnect_0_jtag_uart_pipeline_bridge_s0_byteenable;    // mm_interconnect_0:jtag_uart_pipeline_bridge_s0_byteenable -> jtag_uart_pipeline_bridge:s0_byteenable
	wire         mm_interconnect_0_jtag_uart_pipeline_bridge_s0_readdatavalid; // jtag_uart_pipeline_bridge:s0_readdatavalid -> mm_interconnect_0:jtag_uart_pipeline_bridge_s0_readdatavalid
	wire         mm_interconnect_0_jtag_uart_pipeline_bridge_s0_write;         // mm_interconnect_0:jtag_uart_pipeline_bridge_s0_write -> jtag_uart_pipeline_bridge:s0_write
	wire  [31:0] mm_interconnect_0_jtag_uart_pipeline_bridge_s0_writedata;     // mm_interconnect_0:jtag_uart_pipeline_bridge_s0_writedata -> jtag_uart_pipeline_bridge:s0_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_pipeline_bridge_s0_burstcount;    // mm_interconnect_0:jtag_uart_pipeline_bridge_s0_burstcount -> jtag_uart_pipeline_bridge:s0_burstcount
	wire  [31:0] mm_interconnect_0_pio_pipeline_bridge_s0_readdata;            // pio_pipeline_bridge:s0_readdata -> mm_interconnect_0:pio_pipeline_bridge_s0_readdata
	wire         mm_interconnect_0_pio_pipeline_bridge_s0_waitrequest;         // pio_pipeline_bridge:s0_waitrequest -> mm_interconnect_0:pio_pipeline_bridge_s0_waitrequest
	wire         mm_interconnect_0_pio_pipeline_bridge_s0_debugaccess;         // mm_interconnect_0:pio_pipeline_bridge_s0_debugaccess -> pio_pipeline_bridge:s0_debugaccess
	wire   [3:0] mm_interconnect_0_pio_pipeline_bridge_s0_address;             // mm_interconnect_0:pio_pipeline_bridge_s0_address -> pio_pipeline_bridge:s0_address
	wire         mm_interconnect_0_pio_pipeline_bridge_s0_read;                // mm_interconnect_0:pio_pipeline_bridge_s0_read -> pio_pipeline_bridge:s0_read
	wire   [3:0] mm_interconnect_0_pio_pipeline_bridge_s0_byteenable;          // mm_interconnect_0:pio_pipeline_bridge_s0_byteenable -> pio_pipeline_bridge:s0_byteenable
	wire         mm_interconnect_0_pio_pipeline_bridge_s0_readdatavalid;       // pio_pipeline_bridge:s0_readdatavalid -> mm_interconnect_0:pio_pipeline_bridge_s0_readdatavalid
	wire         mm_interconnect_0_pio_pipeline_bridge_s0_write;               // mm_interconnect_0:pio_pipeline_bridge_s0_write -> pio_pipeline_bridge:s0_write
	wire  [31:0] mm_interconnect_0_pio_pipeline_bridge_s0_writedata;           // mm_interconnect_0:pio_pipeline_bridge_s0_writedata -> pio_pipeline_bridge:s0_writedata
	wire   [0:0] mm_interconnect_0_pio_pipeline_bridge_s0_burstcount;          // mm_interconnect_0:pio_pipeline_bridge_s0_burstcount -> pio_pipeline_bridge:s0_burstcount
	wire         mm_interconnect_0_on_chip_memory_s1_chipselect;               // mm_interconnect_0:on_chip_memory_s1_chipselect -> on_chip_memory:chipselect
	wire  [31:0] mm_interconnect_0_on_chip_memory_s1_readdata;                 // on_chip_memory:readdata -> mm_interconnect_0:on_chip_memory_s1_readdata
	wire   [9:0] mm_interconnect_0_on_chip_memory_s1_address;                  // mm_interconnect_0:on_chip_memory_s1_address -> on_chip_memory:address
	wire   [3:0] mm_interconnect_0_on_chip_memory_s1_byteenable;               // mm_interconnect_0:on_chip_memory_s1_byteenable -> on_chip_memory:byteenable
	wire         mm_interconnect_0_on_chip_memory_s1_write;                    // mm_interconnect_0:on_chip_memory_s1_write -> on_chip_memory:write
	wire  [31:0] mm_interconnect_0_on_chip_memory_s1_writedata;                // mm_interconnect_0:on_chip_memory_s1_writedata -> on_chip_memory:writedata
	wire         mm_interconnect_0_on_chip_memory_s1_clken;                    // mm_interconnect_0:on_chip_memory_s1_clken -> on_chip_memory:clken
	wire         jtag_uart_pipeline_bridge_m0_waitrequest;                     // mm_interconnect_1:jtag_uart_pipeline_bridge_m0_waitrequest -> jtag_uart_pipeline_bridge:m0_waitrequest
	wire  [31:0] jtag_uart_pipeline_bridge_m0_readdata;                        // mm_interconnect_1:jtag_uart_pipeline_bridge_m0_readdata -> jtag_uart_pipeline_bridge:m0_readdata
	wire         jtag_uart_pipeline_bridge_m0_debugaccess;                     // jtag_uart_pipeline_bridge:m0_debugaccess -> mm_interconnect_1:jtag_uart_pipeline_bridge_m0_debugaccess
	wire   [2:0] jtag_uart_pipeline_bridge_m0_address;                         // jtag_uart_pipeline_bridge:m0_address -> mm_interconnect_1:jtag_uart_pipeline_bridge_m0_address
	wire         jtag_uart_pipeline_bridge_m0_read;                            // jtag_uart_pipeline_bridge:m0_read -> mm_interconnect_1:jtag_uart_pipeline_bridge_m0_read
	wire   [3:0] jtag_uart_pipeline_bridge_m0_byteenable;                      // jtag_uart_pipeline_bridge:m0_byteenable -> mm_interconnect_1:jtag_uart_pipeline_bridge_m0_byteenable
	wire         jtag_uart_pipeline_bridge_m0_readdatavalid;                   // mm_interconnect_1:jtag_uart_pipeline_bridge_m0_readdatavalid -> jtag_uart_pipeline_bridge:m0_readdatavalid
	wire  [31:0] jtag_uart_pipeline_bridge_m0_writedata;                       // jtag_uart_pipeline_bridge:m0_writedata -> mm_interconnect_1:jtag_uart_pipeline_bridge_m0_writedata
	wire         jtag_uart_pipeline_bridge_m0_write;                           // jtag_uart_pipeline_bridge:m0_write -> mm_interconnect_1:jtag_uart_pipeline_bridge_m0_write
	wire   [0:0] jtag_uart_pipeline_bridge_m0_burstcount;                      // jtag_uart_pipeline_bridge:m0_burstcount -> mm_interconnect_1:jtag_uart_pipeline_bridge_m0_burstcount
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect;     // mm_interconnect_1:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata;       // jtag_uart:av_readdata -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest;    // jtag_uart:av_waitrequest -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_address;        // mm_interconnect_1:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_read;           // mm_interconnect_1:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_write;          // mm_interconnect_1:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata;      // mm_interconnect_1:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         pio_pipeline_bridge_m0_waitrequest;                           // mm_interconnect_2:pio_pipeline_bridge_m0_waitrequest -> pio_pipeline_bridge:m0_waitrequest
	wire  [31:0] pio_pipeline_bridge_m0_readdata;                              // mm_interconnect_2:pio_pipeline_bridge_m0_readdata -> pio_pipeline_bridge:m0_readdata
	wire         pio_pipeline_bridge_m0_debugaccess;                           // pio_pipeline_bridge:m0_debugaccess -> mm_interconnect_2:pio_pipeline_bridge_m0_debugaccess
	wire   [3:0] pio_pipeline_bridge_m0_address;                               // pio_pipeline_bridge:m0_address -> mm_interconnect_2:pio_pipeline_bridge_m0_address
	wire         pio_pipeline_bridge_m0_read;                                  // pio_pipeline_bridge:m0_read -> mm_interconnect_2:pio_pipeline_bridge_m0_read
	wire   [3:0] pio_pipeline_bridge_m0_byteenable;                            // pio_pipeline_bridge:m0_byteenable -> mm_interconnect_2:pio_pipeline_bridge_m0_byteenable
	wire         pio_pipeline_bridge_m0_readdatavalid;                         // mm_interconnect_2:pio_pipeline_bridge_m0_readdatavalid -> pio_pipeline_bridge:m0_readdatavalid
	wire  [31:0] pio_pipeline_bridge_m0_writedata;                             // pio_pipeline_bridge:m0_writedata -> mm_interconnect_2:pio_pipeline_bridge_m0_writedata
	wire         pio_pipeline_bridge_m0_write;                                 // pio_pipeline_bridge:m0_write -> mm_interconnect_2:pio_pipeline_bridge_m0_write
	wire   [0:0] pio_pipeline_bridge_m0_burstcount;                            // pio_pipeline_bridge:m0_burstcount -> mm_interconnect_2:pio_pipeline_bridge_m0_burstcount
	wire         mm_interconnect_2_leds_s1_chipselect;                         // mm_interconnect_2:leds_s1_chipselect -> leds:chipselect
	wire  [31:0] mm_interconnect_2_leds_s1_readdata;                           // leds:readdata -> mm_interconnect_2:leds_s1_readdata
	wire   [1:0] mm_interconnect_2_leds_s1_address;                            // mm_interconnect_2:leds_s1_address -> leds:address
	wire         mm_interconnect_2_leds_s1_write;                              // mm_interconnect_2:leds_s1_write -> leds:write_n
	wire  [31:0] mm_interconnect_2_leds_s1_writedata;                          // mm_interconnect_2:leds_s1_writedata -> leds:writedata
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [jtag_uart:rst_n, jtag_uart_pipeline_bridge:reset, leds:reset_n, mm_interconnect_0:rv32i_core_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_1:jtag_uart_pipeline_bridge_reset_reset_bridge_in_reset_reset, mm_interconnect_2:pio_pipeline_bridge_reset_reset_bridge_in_reset_reset, on_chip_memory:reset, pio_pipeline_bridge:reset, rst_translator:in_reset, rv32i_core:rst_n]
	wire         rst_controller_reset_out_reset_req;                           // rst_controller:reset_req -> [on_chip_memory:reset_req, rst_translator:reset_req_in]

	soc_simple_PLL_50_150 pll_50_150 (
		.refclk   (clk_clk),                //  refclk.clk
		.rst      (~reset_reset_n),         //   reset.reset
		.outclk_0 (pll_50_150_outclk0_clk), // outclk0.clk
		.locked   (locked_export)           //  locked.export
	);

	soc_simple_jtag_uart jtag_uart (
		.clk            (pll_50_150_outclk0_clk),                                    //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         ()                                                           //               irq.irq
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (3),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) jtag_uart_pipeline_bridge (
		.clk              (pll_50_150_outclk0_clk),                                       //   clk.clk
		.reset            (rst_controller_reset_out_reset),                               // reset.reset
		.s0_waitrequest   (mm_interconnect_0_jtag_uart_pipeline_bridge_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_jtag_uart_pipeline_bridge_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_jtag_uart_pipeline_bridge_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_jtag_uart_pipeline_bridge_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_jtag_uart_pipeline_bridge_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_jtag_uart_pipeline_bridge_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_jtag_uart_pipeline_bridge_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_jtag_uart_pipeline_bridge_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_jtag_uart_pipeline_bridge_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_jtag_uart_pipeline_bridge_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (jtag_uart_pipeline_bridge_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (jtag_uart_pipeline_bridge_m0_readdata),                        //      .readdata
		.m0_readdatavalid (jtag_uart_pipeline_bridge_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (jtag_uart_pipeline_bridge_m0_burstcount),                      //      .burstcount
		.m0_writedata     (jtag_uart_pipeline_bridge_m0_writedata),                       //      .writedata
		.m0_address       (jtag_uart_pipeline_bridge_m0_address),                         //      .address
		.m0_write         (jtag_uart_pipeline_bridge_m0_write),                           //      .write
		.m0_read          (jtag_uart_pipeline_bridge_m0_read),                            //      .read
		.m0_byteenable    (jtag_uart_pipeline_bridge_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (jtag_uart_pipeline_bridge_m0_debugaccess),                     //      .debugaccess
		.s0_response      (),                                                             // (terminated)
		.m0_response      (2'b00)                                                         // (terminated)
	);

	soc_simple_leds leds (
		.clk        (pll_50_150_outclk0_clk),               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_2_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_leds_s1_readdata),   //                    .readdata
		.out_port   (leds_export)                           // external_connection.export
	);

	soc_simple_on_chip_memory on_chip_memory (
		.clk        (pll_50_150_outclk0_clk),                         //   clk1.clk
		.address    (mm_interconnect_0_on_chip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_on_chip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_on_chip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_on_chip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_on_chip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_on_chip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_on_chip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                 // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),             //       .reset_req
		.freeze     (1'b0)                                            // (terminated)
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (4),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) pio_pipeline_bridge (
		.clk              (pll_50_150_outclk0_clk),                                 //   clk.clk
		.reset            (rst_controller_reset_out_reset),                         // reset.reset
		.s0_waitrequest   (mm_interconnect_0_pio_pipeline_bridge_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_pio_pipeline_bridge_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_pio_pipeline_bridge_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_pio_pipeline_bridge_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_pio_pipeline_bridge_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_pio_pipeline_bridge_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_pio_pipeline_bridge_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_pio_pipeline_bridge_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_pio_pipeline_bridge_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_pio_pipeline_bridge_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (pio_pipeline_bridge_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (pio_pipeline_bridge_m0_readdata),                        //      .readdata
		.m0_readdatavalid (pio_pipeline_bridge_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (pio_pipeline_bridge_m0_burstcount),                      //      .burstcount
		.m0_writedata     (pio_pipeline_bridge_m0_writedata),                       //      .writedata
		.m0_address       (pio_pipeline_bridge_m0_address),                         //      .address
		.m0_write         (pio_pipeline_bridge_m0_write),                           //      .write
		.m0_read          (pio_pipeline_bridge_m0_read),                            //      .read
		.m0_byteenable    (pio_pipeline_bridge_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (pio_pipeline_bridge_m0_debugaccess),                     //      .debugaccess
		.s0_response      (),                                                       // (terminated)
		.m0_response      (2'b00)                                                   // (terminated)
	);

	risac_avalon rv32i_core (
		.clk              (pll_50_150_outclk0_clk),                    //              clock.clk
		.rst_n            (~rst_controller_reset_out_reset),           //         reset_sink.reset_n
		.avIB_readdata    (rv32i_core_instruction_master_readdata),    // instruction_master.readdata
		.avIB_address     (rv32i_core_instruction_master_address),     //                   .address
		.avIB_waitrequest (rv32i_core_instruction_master_waitrequest), //                   .waitrequest
		.avIB_read        (rv32i_core_instruction_master_read),        //                   .read
		.avDB_address     (rv32i_core_data_master_address),            //        data_master.address
		.avDB_readdata    (rv32i_core_data_master_readdata),           //                   .readdata
		.avDB_read        (rv32i_core_data_master_read),               //                   .read
		.avDB_writedata   (rv32i_core_data_master_writedata),          //                   .writedata
		.avDB_byteenable  (rv32i_core_data_master_byteenable),         //                   .byteenable
		.avDB_write       (rv32i_core_data_master_write),              //                   .write
		.avDB_waitrequest (rv32i_core_data_master_waitrequest)         //                   .waitrequest
	);

	soc_simple_mm_interconnect_0 mm_interconnect_0 (
		.PLL_50_150_outclk0_clk                            (pll_50_150_outclk0_clk),                                       //                          PLL_50_150_outclk0.clk
		.rv32i_core_reset_sink_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                               // rv32i_core_reset_sink_reset_bridge_in_reset.reset
		.rv32i_core_data_master_address                    (rv32i_core_data_master_address),                               //                      rv32i_core_data_master.address
		.rv32i_core_data_master_waitrequest                (rv32i_core_data_master_waitrequest),                           //                                            .waitrequest
		.rv32i_core_data_master_byteenable                 (rv32i_core_data_master_byteenable),                            //                                            .byteenable
		.rv32i_core_data_master_read                       (rv32i_core_data_master_read),                                  //                                            .read
		.rv32i_core_data_master_readdata                   (rv32i_core_data_master_readdata),                              //                                            .readdata
		.rv32i_core_data_master_write                      (rv32i_core_data_master_write),                                 //                                            .write
		.rv32i_core_data_master_writedata                  (rv32i_core_data_master_writedata),                             //                                            .writedata
		.rv32i_core_instruction_master_address             (rv32i_core_instruction_master_address),                        //               rv32i_core_instruction_master.address
		.rv32i_core_instruction_master_waitrequest         (rv32i_core_instruction_master_waitrequest),                    //                                            .waitrequest
		.rv32i_core_instruction_master_read                (rv32i_core_instruction_master_read),                           //                                            .read
		.rv32i_core_instruction_master_readdata            (rv32i_core_instruction_master_readdata),                       //                                            .readdata
		.jtag_uart_pipeline_bridge_s0_address              (mm_interconnect_0_jtag_uart_pipeline_bridge_s0_address),       //                jtag_uart_pipeline_bridge_s0.address
		.jtag_uart_pipeline_bridge_s0_write                (mm_interconnect_0_jtag_uart_pipeline_bridge_s0_write),         //                                            .write
		.jtag_uart_pipeline_bridge_s0_read                 (mm_interconnect_0_jtag_uart_pipeline_bridge_s0_read),          //                                            .read
		.jtag_uart_pipeline_bridge_s0_readdata             (mm_interconnect_0_jtag_uart_pipeline_bridge_s0_readdata),      //                                            .readdata
		.jtag_uart_pipeline_bridge_s0_writedata            (mm_interconnect_0_jtag_uart_pipeline_bridge_s0_writedata),     //                                            .writedata
		.jtag_uart_pipeline_bridge_s0_burstcount           (mm_interconnect_0_jtag_uart_pipeline_bridge_s0_burstcount),    //                                            .burstcount
		.jtag_uart_pipeline_bridge_s0_byteenable           (mm_interconnect_0_jtag_uart_pipeline_bridge_s0_byteenable),    //                                            .byteenable
		.jtag_uart_pipeline_bridge_s0_readdatavalid        (mm_interconnect_0_jtag_uart_pipeline_bridge_s0_readdatavalid), //                                            .readdatavalid
		.jtag_uart_pipeline_bridge_s0_waitrequest          (mm_interconnect_0_jtag_uart_pipeline_bridge_s0_waitrequest),   //                                            .waitrequest
		.jtag_uart_pipeline_bridge_s0_debugaccess          (mm_interconnect_0_jtag_uart_pipeline_bridge_s0_debugaccess),   //                                            .debugaccess
		.on_chip_memory_s1_address                         (mm_interconnect_0_on_chip_memory_s1_address),                  //                           on_chip_memory_s1.address
		.on_chip_memory_s1_write                           (mm_interconnect_0_on_chip_memory_s1_write),                    //                                            .write
		.on_chip_memory_s1_readdata                        (mm_interconnect_0_on_chip_memory_s1_readdata),                 //                                            .readdata
		.on_chip_memory_s1_writedata                       (mm_interconnect_0_on_chip_memory_s1_writedata),                //                                            .writedata
		.on_chip_memory_s1_byteenable                      (mm_interconnect_0_on_chip_memory_s1_byteenable),               //                                            .byteenable
		.on_chip_memory_s1_chipselect                      (mm_interconnect_0_on_chip_memory_s1_chipselect),               //                                            .chipselect
		.on_chip_memory_s1_clken                           (mm_interconnect_0_on_chip_memory_s1_clken),                    //                                            .clken
		.pio_pipeline_bridge_s0_address                    (mm_interconnect_0_pio_pipeline_bridge_s0_address),             //                      pio_pipeline_bridge_s0.address
		.pio_pipeline_bridge_s0_write                      (mm_interconnect_0_pio_pipeline_bridge_s0_write),               //                                            .write
		.pio_pipeline_bridge_s0_read                       (mm_interconnect_0_pio_pipeline_bridge_s0_read),                //                                            .read
		.pio_pipeline_bridge_s0_readdata                   (mm_interconnect_0_pio_pipeline_bridge_s0_readdata),            //                                            .readdata
		.pio_pipeline_bridge_s0_writedata                  (mm_interconnect_0_pio_pipeline_bridge_s0_writedata),           //                                            .writedata
		.pio_pipeline_bridge_s0_burstcount                 (mm_interconnect_0_pio_pipeline_bridge_s0_burstcount),          //                                            .burstcount
		.pio_pipeline_bridge_s0_byteenable                 (mm_interconnect_0_pio_pipeline_bridge_s0_byteenable),          //                                            .byteenable
		.pio_pipeline_bridge_s0_readdatavalid              (mm_interconnect_0_pio_pipeline_bridge_s0_readdatavalid),       //                                            .readdatavalid
		.pio_pipeline_bridge_s0_waitrequest                (mm_interconnect_0_pio_pipeline_bridge_s0_waitrequest),         //                                            .waitrequest
		.pio_pipeline_bridge_s0_debugaccess                (mm_interconnect_0_pio_pipeline_bridge_s0_debugaccess)          //                                            .debugaccess
	);

	soc_simple_mm_interconnect_1 mm_interconnect_1 (
		.PLL_50_150_outclk0_clk                                      (pll_50_150_outclk0_clk),                                    //                                    PLL_50_150_outclk0.clk
		.jtag_uart_pipeline_bridge_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // jtag_uart_pipeline_bridge_reset_reset_bridge_in_reset.reset
		.jtag_uart_pipeline_bridge_m0_address                        (jtag_uart_pipeline_bridge_m0_address),                      //                          jtag_uart_pipeline_bridge_m0.address
		.jtag_uart_pipeline_bridge_m0_waitrequest                    (jtag_uart_pipeline_bridge_m0_waitrequest),                  //                                                      .waitrequest
		.jtag_uart_pipeline_bridge_m0_burstcount                     (jtag_uart_pipeline_bridge_m0_burstcount),                   //                                                      .burstcount
		.jtag_uart_pipeline_bridge_m0_byteenable                     (jtag_uart_pipeline_bridge_m0_byteenable),                   //                                                      .byteenable
		.jtag_uart_pipeline_bridge_m0_read                           (jtag_uart_pipeline_bridge_m0_read),                         //                                                      .read
		.jtag_uart_pipeline_bridge_m0_readdata                       (jtag_uart_pipeline_bridge_m0_readdata),                     //                                                      .readdata
		.jtag_uart_pipeline_bridge_m0_readdatavalid                  (jtag_uart_pipeline_bridge_m0_readdatavalid),                //                                                      .readdatavalid
		.jtag_uart_pipeline_bridge_m0_write                          (jtag_uart_pipeline_bridge_m0_write),                        //                                                      .write
		.jtag_uart_pipeline_bridge_m0_writedata                      (jtag_uart_pipeline_bridge_m0_writedata),                    //                                                      .writedata
		.jtag_uart_pipeline_bridge_m0_debugaccess                    (jtag_uart_pipeline_bridge_m0_debugaccess),                  //                                                      .debugaccess
		.jtag_uart_avalon_jtag_slave_address                         (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                           jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                           (mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),       //                                                      .write
		.jtag_uart_avalon_jtag_slave_read                            (mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),        //                                                      .read
		.jtag_uart_avalon_jtag_slave_readdata                        (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                                                      .readdata
		.jtag_uart_avalon_jtag_slave_writedata                       (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                                                      .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                                                      .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                      (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect)   //                                                      .chipselect
	);

	soc_simple_mm_interconnect_2 mm_interconnect_2 (
		.PLL_50_150_outclk0_clk                                (pll_50_150_outclk0_clk),               //                              PLL_50_150_outclk0.clk
		.pio_pipeline_bridge_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),       // pio_pipeline_bridge_reset_reset_bridge_in_reset.reset
		.pio_pipeline_bridge_m0_address                        (pio_pipeline_bridge_m0_address),       //                          pio_pipeline_bridge_m0.address
		.pio_pipeline_bridge_m0_waitrequest                    (pio_pipeline_bridge_m0_waitrequest),   //                                                .waitrequest
		.pio_pipeline_bridge_m0_burstcount                     (pio_pipeline_bridge_m0_burstcount),    //                                                .burstcount
		.pio_pipeline_bridge_m0_byteenable                     (pio_pipeline_bridge_m0_byteenable),    //                                                .byteenable
		.pio_pipeline_bridge_m0_read                           (pio_pipeline_bridge_m0_read),          //                                                .read
		.pio_pipeline_bridge_m0_readdata                       (pio_pipeline_bridge_m0_readdata),      //                                                .readdata
		.pio_pipeline_bridge_m0_readdatavalid                  (pio_pipeline_bridge_m0_readdatavalid), //                                                .readdatavalid
		.pio_pipeline_bridge_m0_write                          (pio_pipeline_bridge_m0_write),         //                                                .write
		.pio_pipeline_bridge_m0_writedata                      (pio_pipeline_bridge_m0_writedata),     //                                                .writedata
		.pio_pipeline_bridge_m0_debugaccess                    (pio_pipeline_bridge_m0_debugaccess),   //                                                .debugaccess
		.leds_s1_address                                       (mm_interconnect_2_leds_s1_address),    //                                         leds_s1.address
		.leds_s1_write                                         (mm_interconnect_2_leds_s1_write),      //                                                .write
		.leds_s1_readdata                                      (mm_interconnect_2_leds_s1_readdata),   //                                                .readdata
		.leds_s1_writedata                                     (mm_interconnect_2_leds_s1_writedata),  //                                                .writedata
		.leds_s1_chipselect                                    (mm_interconnect_2_leds_s1_chipselect)  //                                                .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (pll_50_150_outclk0_clk),             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
