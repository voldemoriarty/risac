// risac_soc_system.v

// Generated using ACDS version 13.0 156 at 2019.11.15.16:54:40

`timescale 1 ps / 1 ps
module risac_soc_system (
		input  wire       clk_clk,       //   clk.clk
		input  wire       reset_reset_n, // reset.reset_n
		output wire [9:0] ledr_export,   //  ledr.export
		input  wire       uart_rxd,      //  uart.rxd
		output wire       uart_txd       //      .txd
	);

	wire          rv32i_core_instruction_master_waitrequest;                                                 // RV32I_Core_instruction_master_translator:av_waitrequest -> RV32I_Core:avIB_waitrequest
	wire   [31:0] rv32i_core_instruction_master_address;                                                     // RV32I_Core:avIB_address -> RV32I_Core_instruction_master_translator:av_address
	wire          rv32i_core_instruction_master_read;                                                        // RV32I_Core:avIB_read -> RV32I_Core_instruction_master_translator:av_read
	wire   [31:0] rv32i_core_instruction_master_readdata;                                                    // RV32I_Core_instruction_master_translator:av_readdata -> RV32I_Core:avIB_readdata
	wire          rv32i_core_data_master_waitrequest;                                                        // RV32I_Core_data_master_translator:av_waitrequest -> RV32I_Core:avDB_waitrequest
	wire   [31:0] rv32i_core_data_master_writedata;                                                          // RV32I_Core:avDB_writedata -> RV32I_Core_data_master_translator:av_writedata
	wire   [31:0] rv32i_core_data_master_address;                                                            // RV32I_Core:avDB_address -> RV32I_Core_data_master_translator:av_address
	wire          rv32i_core_data_master_write;                                                              // RV32I_Core:avDB_write -> RV32I_Core_data_master_translator:av_write
	wire          rv32i_core_data_master_read;                                                               // RV32I_Core:avDB_read -> RV32I_Core_data_master_translator:av_read
	wire   [31:0] rv32i_core_data_master_readdata;                                                           // RV32I_Core_data_master_translator:av_readdata -> RV32I_Core:avDB_readdata
	wire    [3:0] rv32i_core_data_master_byteenable;                                                         // RV32I_Core:avDB_byteenable -> RV32I_Core_data_master_translator:av_byteenable
	wire   [31:0] memory_s1_translator_avalon_anti_slave_0_writedata;                                        // Memory_s1_translator:av_writedata -> Memory:writedata
	wire    [9:0] memory_s1_translator_avalon_anti_slave_0_address;                                          // Memory_s1_translator:av_address -> Memory:address
	wire          memory_s1_translator_avalon_anti_slave_0_chipselect;                                       // Memory_s1_translator:av_chipselect -> Memory:chipselect
	wire          memory_s1_translator_avalon_anti_slave_0_clken;                                            // Memory_s1_translator:av_clken -> Memory:clken
	wire          memory_s1_translator_avalon_anti_slave_0_write;                                            // Memory_s1_translator:av_write -> Memory:write
	wire   [31:0] memory_s1_translator_avalon_anti_slave_0_readdata;                                         // Memory:readdata -> Memory_s1_translator:av_readdata
	wire    [3:0] memory_s1_translator_avalon_anti_slave_0_byteenable;                                       // Memory_s1_translator:av_byteenable -> Memory:byteenable
	wire   [31:0] ledr_s1_translator_avalon_anti_slave_0_writedata;                                          // LEDR_s1_translator:av_writedata -> LEDR:writedata
	wire    [1:0] ledr_s1_translator_avalon_anti_slave_0_address;                                            // LEDR_s1_translator:av_address -> LEDR:address
	wire          ledr_s1_translator_avalon_anti_slave_0_chipselect;                                         // LEDR_s1_translator:av_chipselect -> LEDR:chipselect
	wire          ledr_s1_translator_avalon_anti_slave_0_write;                                              // LEDR_s1_translator:av_write -> LEDR:write_n
	wire   [31:0] ledr_s1_translator_avalon_anti_slave_0_readdata;                                           // LEDR:readdata -> LEDR_s1_translator:av_readdata
	wire   [15:0] uart_0_s1_translator_avalon_anti_slave_0_writedata;                                        // uart_0_s1_translator:av_writedata -> uart_0:writedata
	wire    [2:0] uart_0_s1_translator_avalon_anti_slave_0_address;                                          // uart_0_s1_translator:av_address -> uart_0:address
	wire          uart_0_s1_translator_avalon_anti_slave_0_chipselect;                                       // uart_0_s1_translator:av_chipselect -> uart_0:chipselect
	wire          uart_0_s1_translator_avalon_anti_slave_0_write;                                            // uart_0_s1_translator:av_write -> uart_0:write_n
	wire          uart_0_s1_translator_avalon_anti_slave_0_read;                                             // uart_0_s1_translator:av_read -> uart_0:read_n
	wire   [15:0] uart_0_s1_translator_avalon_anti_slave_0_readdata;                                         // uart_0:readdata -> uart_0_s1_translator:av_readdata
	wire          uart_0_s1_translator_avalon_anti_slave_0_begintransfer;                                    // uart_0_s1_translator:av_begintransfer -> uart_0:begintransfer
	wire          rv32i_core_instruction_master_translator_avalon_universal_master_0_waitrequest;            // RV32I_Core_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> RV32I_Core_instruction_master_translator:uav_waitrequest
	wire    [2:0] rv32i_core_instruction_master_translator_avalon_universal_master_0_burstcount;             // RV32I_Core_instruction_master_translator:uav_burstcount -> RV32I_Core_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] rv32i_core_instruction_master_translator_avalon_universal_master_0_writedata;              // RV32I_Core_instruction_master_translator:uav_writedata -> RV32I_Core_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] rv32i_core_instruction_master_translator_avalon_universal_master_0_address;                // RV32I_Core_instruction_master_translator:uav_address -> RV32I_Core_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          rv32i_core_instruction_master_translator_avalon_universal_master_0_lock;                   // RV32I_Core_instruction_master_translator:uav_lock -> RV32I_Core_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          rv32i_core_instruction_master_translator_avalon_universal_master_0_write;                  // RV32I_Core_instruction_master_translator:uav_write -> RV32I_Core_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          rv32i_core_instruction_master_translator_avalon_universal_master_0_read;                   // RV32I_Core_instruction_master_translator:uav_read -> RV32I_Core_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] rv32i_core_instruction_master_translator_avalon_universal_master_0_readdata;               // RV32I_Core_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> RV32I_Core_instruction_master_translator:uav_readdata
	wire          rv32i_core_instruction_master_translator_avalon_universal_master_0_debugaccess;            // RV32I_Core_instruction_master_translator:uav_debugaccess -> RV32I_Core_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] rv32i_core_instruction_master_translator_avalon_universal_master_0_byteenable;             // RV32I_Core_instruction_master_translator:uav_byteenable -> RV32I_Core_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          rv32i_core_instruction_master_translator_avalon_universal_master_0_readdatavalid;          // RV32I_Core_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> RV32I_Core_instruction_master_translator:uav_readdatavalid
	wire          rv32i_core_data_master_translator_avalon_universal_master_0_waitrequest;                   // RV32I_Core_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> RV32I_Core_data_master_translator:uav_waitrequest
	wire    [2:0] rv32i_core_data_master_translator_avalon_universal_master_0_burstcount;                    // RV32I_Core_data_master_translator:uav_burstcount -> RV32I_Core_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] rv32i_core_data_master_translator_avalon_universal_master_0_writedata;                     // RV32I_Core_data_master_translator:uav_writedata -> RV32I_Core_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] rv32i_core_data_master_translator_avalon_universal_master_0_address;                       // RV32I_Core_data_master_translator:uav_address -> RV32I_Core_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          rv32i_core_data_master_translator_avalon_universal_master_0_lock;                          // RV32I_Core_data_master_translator:uav_lock -> RV32I_Core_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          rv32i_core_data_master_translator_avalon_universal_master_0_write;                         // RV32I_Core_data_master_translator:uav_write -> RV32I_Core_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          rv32i_core_data_master_translator_avalon_universal_master_0_read;                          // RV32I_Core_data_master_translator:uav_read -> RV32I_Core_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] rv32i_core_data_master_translator_avalon_universal_master_0_readdata;                      // RV32I_Core_data_master_translator_avalon_universal_master_0_agent:av_readdata -> RV32I_Core_data_master_translator:uav_readdata
	wire          rv32i_core_data_master_translator_avalon_universal_master_0_debugaccess;                   // RV32I_Core_data_master_translator:uav_debugaccess -> RV32I_Core_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] rv32i_core_data_master_translator_avalon_universal_master_0_byteenable;                    // RV32I_Core_data_master_translator:uav_byteenable -> RV32I_Core_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          rv32i_core_data_master_translator_avalon_universal_master_0_readdatavalid;                 // RV32I_Core_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> RV32I_Core_data_master_translator:uav_readdatavalid
	wire          memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // Memory_s1_translator:uav_waitrequest -> Memory_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // Memory_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> Memory_s1_translator:uav_burstcount
	wire   [31:0] memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                          // Memory_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> Memory_s1_translator:uav_writedata
	wire   [31:0] memory_s1_translator_avalon_universal_slave_0_agent_m0_address;                            // Memory_s1_translator_avalon_universal_slave_0_agent:m0_address -> Memory_s1_translator:uav_address
	wire          memory_s1_translator_avalon_universal_slave_0_agent_m0_write;                              // Memory_s1_translator_avalon_universal_slave_0_agent:m0_write -> Memory_s1_translator:uav_write
	wire          memory_s1_translator_avalon_universal_slave_0_agent_m0_lock;                               // Memory_s1_translator_avalon_universal_slave_0_agent:m0_lock -> Memory_s1_translator:uav_lock
	wire          memory_s1_translator_avalon_universal_slave_0_agent_m0_read;                               // Memory_s1_translator_avalon_universal_slave_0_agent:m0_read -> Memory_s1_translator:uav_read
	wire   [31:0] memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                           // Memory_s1_translator:uav_readdata -> Memory_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // Memory_s1_translator:uav_readdatavalid -> Memory_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // Memory_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Memory_s1_translator:uav_debugaccess
	wire    [3:0] memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // Memory_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> Memory_s1_translator:uav_byteenable
	wire          memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // Memory_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // Memory_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // Memory_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [101:0] memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                        // Memory_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Memory_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [101:0] memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // Memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // Memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // Memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // Memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                          // LEDR_s1_translator:uav_waitrequest -> LEDR_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                           // LEDR_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> LEDR_s1_translator:uav_burstcount
	wire   [31:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                            // LEDR_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> LEDR_s1_translator:uav_writedata
	wire   [31:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_address;                              // LEDR_s1_translator_avalon_universal_slave_0_agent:m0_address -> LEDR_s1_translator:uav_address
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_m0_write;                                // LEDR_s1_translator_avalon_universal_slave_0_agent:m0_write -> LEDR_s1_translator:uav_write
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                 // LEDR_s1_translator_avalon_universal_slave_0_agent:m0_lock -> LEDR_s1_translator:uav_lock
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_m0_read;                                 // LEDR_s1_translator_avalon_universal_slave_0_agent:m0_read -> LEDR_s1_translator:uav_read
	wire   [31:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                             // LEDR_s1_translator:uav_readdata -> LEDR_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                        // LEDR_s1_translator:uav_readdatavalid -> LEDR_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                          // LEDR_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> LEDR_s1_translator:uav_debugaccess
	wire    [3:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                           // LEDR_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> LEDR_s1_translator:uav_byteenable
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                   // LEDR_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                         // LEDR_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                 // LEDR_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [101:0] ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                          // LEDR_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                         // LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> LEDR_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                // LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> LEDR_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                      // LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> LEDR_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;              // LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> LEDR_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [101:0] ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                       // LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> LEDR_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                      // LEDR_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                    // LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                     // LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                    // LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // uart_0_s1_translator:uav_waitrequest -> uart_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] uart_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> uart_0_s1_translator:uav_burstcount
	wire   [31:0] uart_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                          // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> uart_0_s1_translator:uav_writedata
	wire   [31:0] uart_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                            // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> uart_0_s1_translator:uav_address
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                              // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> uart_0_s1_translator:uav_write
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                               // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> uart_0_s1_translator:uav_lock
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                               // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> uart_0_s1_translator:uav_read
	wire   [31:0] uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                           // uart_0_s1_translator:uav_readdata -> uart_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // uart_0_s1_translator:uav_readdatavalid -> uart_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> uart_0_s1_translator:uav_debugaccess
	wire    [3:0] uart_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> uart_0_s1_translator:uav_byteenable
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [101:0] uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                        // uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [101:0] uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          rv32i_core_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;   // RV32I_Core_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          rv32i_core_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;         // RV32I_Core_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          rv32i_core_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket; // RV32I_Core_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [100:0] rv32i_core_instruction_master_translator_avalon_universal_master_0_agent_cp_data;          // RV32I_Core_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          rv32i_core_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;         // addr_router:sink_ready -> RV32I_Core_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          rv32i_core_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;          // RV32I_Core_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          rv32i_core_data_master_translator_avalon_universal_master_0_agent_cp_valid;                // RV32I_Core_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          rv32i_core_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;        // RV32I_Core_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [100:0] rv32i_core_data_master_translator_avalon_universal_master_0_agent_cp_data;                 // RV32I_Core_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          rv32i_core_data_master_translator_avalon_universal_master_0_agent_cp_ready;                // addr_router_001:sink_ready -> RV32I_Core_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // Memory_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          memory_s1_translator_avalon_universal_slave_0_agent_rp_valid;                              // Memory_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // Memory_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [100:0] memory_s1_translator_avalon_universal_slave_0_agent_rp_data;                               // Memory_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          memory_s1_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router:sink_ready -> Memory_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                          // LEDR_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                // LEDR_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                        // LEDR_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [100:0] ledr_s1_translator_avalon_universal_slave_0_agent_rp_data;                                 // LEDR_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          ledr_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                // id_router_001:sink_ready -> LEDR_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // uart_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                              // uart_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // uart_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [100:0] uart_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                               // uart_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_002:sink_ready -> uart_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          rst_controller_reset_out_reset;                                                            // rst_controller:reset_out -> [LEDR:reset_n, LEDR_s1_translator:reset, LEDR_s1_translator_avalon_universal_slave_0_agent:reset, LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Memory:reset, Memory_s1_translator:reset, Memory_s1_translator_avalon_universal_slave_0_agent:reset, Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, RV32I_Core:rst_n, RV32I_Core_data_master_translator:reset, RV32I_Core_data_master_translator_avalon_universal_master_0_agent:reset, RV32I_Core_instruction_master_translator:reset, RV32I_Core_instruction_master_translator_avalon_universal_master_0_agent:reset, addr_router:reset, addr_router_001:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, id_router:reset, id_router_001:reset, id_router_002:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_mux_001:reset, uart_0:reset_n, uart_0_s1_translator:reset, uart_0_s1_translator_avalon_universal_slave_0_agent:reset, uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire          cmd_xbar_demux_src0_endofpacket;                                                           // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                 // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                         // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [100:0] cmd_xbar_demux_src0_data;                                                                  // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire    [2:0] cmd_xbar_demux_src0_channel;                                                               // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire          cmd_xbar_demux_src0_ready;                                                                 // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                       // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                             // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                     // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [100:0] cmd_xbar_demux_001_src0_data;                                                              // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire    [2:0] cmd_xbar_demux_001_src0_channel;                                                           // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                             // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_001_src1_endofpacket;                                                       // cmd_xbar_demux_001:src1_endofpacket -> LEDR_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src1_valid;                                                             // cmd_xbar_demux_001:src1_valid -> LEDR_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src1_startofpacket;                                                     // cmd_xbar_demux_001:src1_startofpacket -> LEDR_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [100:0] cmd_xbar_demux_001_src1_data;                                                              // cmd_xbar_demux_001:src1_data -> LEDR_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [2:0] cmd_xbar_demux_001_src1_channel;                                                           // cmd_xbar_demux_001:src1_channel -> LEDR_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src2_endofpacket;                                                       // cmd_xbar_demux_001:src2_endofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src2_valid;                                                             // cmd_xbar_demux_001:src2_valid -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src2_startofpacket;                                                     // cmd_xbar_demux_001:src2_startofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [100:0] cmd_xbar_demux_001_src2_data;                                                              // cmd_xbar_demux_001:src2_data -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [2:0] cmd_xbar_demux_001_src2_channel;                                                           // cmd_xbar_demux_001:src2_channel -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rsp_xbar_demux_src0_endofpacket;                                                           // rsp_xbar_demux:src0_endofpacket -> RV32I_Core_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                 // rsp_xbar_demux:src0_valid -> RV32I_Core_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                         // rsp_xbar_demux:src0_startofpacket -> RV32I_Core_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [100:0] rsp_xbar_demux_src0_data;                                                                  // rsp_xbar_demux:src0_data -> RV32I_Core_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [2:0] rsp_xbar_demux_src0_channel;                                                               // rsp_xbar_demux:src0_channel -> RV32I_Core_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_src1_endofpacket;                                                           // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                                 // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                                         // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [100:0] rsp_xbar_demux_src1_data;                                                                  // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire    [2:0] rsp_xbar_demux_src1_channel;                                                               // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire          rsp_xbar_demux_src1_ready;                                                                 // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                       // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                             // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux_001:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                     // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [100:0] rsp_xbar_demux_001_src0_data;                                                              // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux_001:sink1_data
	wire    [2:0] rsp_xbar_demux_001_src0_channel;                                                           // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux_001:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                             // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                       // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                             // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux_001:sink2_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                     // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [100:0] rsp_xbar_demux_002_src0_data;                                                              // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux_001:sink2_data
	wire    [2:0] rsp_xbar_demux_002_src0_channel;                                                           // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux_001:sink2_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                             // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire          addr_router_src_endofpacket;                                                               // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          addr_router_src_valid;                                                                     // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire          addr_router_src_startofpacket;                                                             // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [100:0] addr_router_src_data;                                                                      // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire    [2:0] addr_router_src_channel;                                                                   // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire          addr_router_src_ready;                                                                     // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire          rsp_xbar_demux_src0_ready;                                                                 // RV32I_Core_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux:src0_ready
	wire          addr_router_001_src_endofpacket;                                                           // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          addr_router_001_src_valid;                                                                 // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire          addr_router_001_src_startofpacket;                                                         // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [100:0] addr_router_001_src_data;                                                                  // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire    [2:0] addr_router_001_src_channel;                                                               // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire          addr_router_001_src_ready;                                                                 // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire          rsp_xbar_mux_001_src_endofpacket;                                                          // rsp_xbar_mux_001:src_endofpacket -> RV32I_Core_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_001_src_valid;                                                                // rsp_xbar_mux_001:src_valid -> RV32I_Core_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_001_src_startofpacket;                                                        // rsp_xbar_mux_001:src_startofpacket -> RV32I_Core_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [100:0] rsp_xbar_mux_001_src_data;                                                                 // rsp_xbar_mux_001:src_data -> RV32I_Core_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [2:0] rsp_xbar_mux_001_src_channel;                                                              // rsp_xbar_mux_001:src_channel -> RV32I_Core_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_001_src_ready;                                                                // RV32I_Core_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	wire          cmd_xbar_mux_src_endofpacket;                                                              // cmd_xbar_mux:src_endofpacket -> Memory_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                                    // cmd_xbar_mux:src_valid -> Memory_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                            // cmd_xbar_mux:src_startofpacket -> Memory_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [100:0] cmd_xbar_mux_src_data;                                                                     // cmd_xbar_mux:src_data -> Memory_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [2:0] cmd_xbar_mux_src_channel;                                                                  // cmd_xbar_mux:src_channel -> Memory_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_src_ready;                                                                    // Memory_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire          id_router_src_endofpacket;                                                                 // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                       // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                               // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [100:0] id_router_src_data;                                                                        // id_router:src_data -> rsp_xbar_demux:sink_data
	wire    [2:0] id_router_src_channel;                                                                     // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                       // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_demux_001_src1_ready;                                                             // LEDR_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src1_ready
	wire          id_router_001_src_endofpacket;                                                             // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          id_router_001_src_valid;                                                                   // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire          id_router_001_src_startofpacket;                                                           // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [100:0] id_router_001_src_data;                                                                    // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire    [2:0] id_router_001_src_channel;                                                                 // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire          id_router_001_src_ready;                                                                   // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire          cmd_xbar_demux_001_src2_ready;                                                             // uart_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src2_ready
	wire          id_router_002_src_endofpacket;                                                             // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                   // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                           // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [100:0] id_router_002_src_data;                                                                    // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire    [2:0] id_router_002_src_channel;                                                                 // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                   // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready

	risac_avalon rv32i_core (
		.clk              (clk_clk),                                   //              clock.clk
		.rst_n            (~rst_controller_reset_out_reset),           //         reset_sink.reset_n
		.avIB_readdata    (rv32i_core_instruction_master_readdata),    // instruction_master.readdata
		.avIB_address     (rv32i_core_instruction_master_address),     //                   .address
		.avIB_waitrequest (rv32i_core_instruction_master_waitrequest), //                   .waitrequest
		.avIB_read        (rv32i_core_instruction_master_read),        //                   .read
		.avDB_address     (rv32i_core_data_master_address),            //        data_master.address
		.avDB_readdata    (rv32i_core_data_master_readdata),           //                   .readdata
		.avDB_read        (rv32i_core_data_master_read),               //                   .read
		.avDB_writedata   (rv32i_core_data_master_writedata),          //                   .writedata
		.avDB_byteenable  (rv32i_core_data_master_byteenable),         //                   .byteenable
		.avDB_write       (rv32i_core_data_master_write),              //                   .write
		.avDB_waitrequest (rv32i_core_data_master_waitrequest)         //                   .waitrequest
	);

	risac_soc_system_Memory memory (
		.clk        (clk_clk),                                             //   clk1.clk
		.address    (memory_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.clken      (memory_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.chipselect (memory_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.write      (memory_s1_translator_avalon_anti_slave_0_write),      //       .write
		.readdata   (memory_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.writedata  (memory_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (memory_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset)                       // reset1.reset
	);

	risac_soc_system_LEDR ledr (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (ledr_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ledr_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ledr_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ledr_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ledr_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (ledr_export)                                        // external_connection.export
	);

	risac_soc_system_uart_0 uart_0 (
		.clk           (clk_clk),                                                //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                        //               reset.reset_n
		.address       (uart_0_s1_translator_avalon_anti_slave_0_address),       //                  s1.address
		.begintransfer (uart_0_s1_translator_avalon_anti_slave_0_begintransfer), //                    .begintransfer
		.chipselect    (uart_0_s1_translator_avalon_anti_slave_0_chipselect),    //                    .chipselect
		.read_n        (~uart_0_s1_translator_avalon_anti_slave_0_read),         //                    .read_n
		.write_n       (~uart_0_s1_translator_avalon_anti_slave_0_write),        //                    .write_n
		.writedata     (uart_0_s1_translator_avalon_anti_slave_0_writedata),     //                    .writedata
		.readdata      (uart_0_s1_translator_avalon_anti_slave_0_readdata),      //                    .readdata
		.dataavailable (),                                                       //                    .dataavailable
		.readyfordata  (),                                                       //                    .readyfordata
		.rxd           (uart_rxd),                                               // external_connection.export
		.txd           (uart_txd),                                               //                    .export
		.irq           ()                                                        //                 irq.irq
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) rv32i_core_instruction_master_translator (
		.clk                      (clk_clk),                                                                          //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                   //                     reset.reset
		.uav_address              (rv32i_core_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (rv32i_core_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (rv32i_core_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (rv32i_core_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (rv32i_core_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (rv32i_core_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (rv32i_core_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (rv32i_core_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (rv32i_core_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (rv32i_core_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (rv32i_core_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (rv32i_core_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (rv32i_core_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (rv32i_core_instruction_master_read),                                               //                          .read
		.av_readdata              (rv32i_core_instruction_master_readdata),                                           //                          .readdata
		.av_burstcount            (1'b1),                                                                             //               (terminated)
		.av_byteenable            (4'b1111),                                                                          //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                             //               (terminated)
		.av_begintransfer         (1'b0),                                                                             //               (terminated)
		.av_chipselect            (1'b0),                                                                             //               (terminated)
		.av_readdatavalid         (),                                                                                 //               (terminated)
		.av_write                 (1'b0),                                                                             //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                             //               (terminated)
		.av_lock                  (1'b0),                                                                             //               (terminated)
		.av_debugaccess           (1'b0),                                                                             //               (terminated)
		.uav_clken                (),                                                                                 //               (terminated)
		.av_clken                 (1'b1),                                                                             //               (terminated)
		.uav_response             (2'b00),                                                                            //               (terminated)
		.av_response              (),                                                                                 //               (terminated)
		.uav_writeresponserequest (),                                                                                 //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                             //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                             //               (terminated)
		.av_writeresponsevalid    ()                                                                                  //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) rv32i_core_data_master_translator (
		.clk                      (clk_clk),                                                                   //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                            //                     reset.reset
		.uav_address              (rv32i_core_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (rv32i_core_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (rv32i_core_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (rv32i_core_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (rv32i_core_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (rv32i_core_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (rv32i_core_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (rv32i_core_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (rv32i_core_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (rv32i_core_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (rv32i_core_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (rv32i_core_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (rv32i_core_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (rv32i_core_data_master_byteenable),                                         //                          .byteenable
		.av_read                  (rv32i_core_data_master_read),                                               //                          .read
		.av_readdata              (rv32i_core_data_master_readdata),                                           //                          .readdata
		.av_write                 (rv32i_core_data_master_write),                                              //                          .write
		.av_writedata             (rv32i_core_data_master_writedata),                                          //                          .writedata
		.av_burstcount            (1'b1),                                                                      //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                      //               (terminated)
		.av_begintransfer         (1'b0),                                                                      //               (terminated)
		.av_chipselect            (1'b0),                                                                      //               (terminated)
		.av_readdatavalid         (),                                                                          //               (terminated)
		.av_lock                  (1'b0),                                                                      //               (terminated)
		.av_debugaccess           (1'b0),                                                                      //               (terminated)
		.uav_clken                (),                                                                          //               (terminated)
		.av_clken                 (1'b1),                                                                      //               (terminated)
		.uav_response             (2'b00),                                                                     //               (terminated)
		.av_response              (),                                                                          //               (terminated)
		.uav_writeresponserequest (),                                                                          //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                      //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                      //               (terminated)
		.av_writeresponsevalid    ()                                                                           //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (10),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) memory_s1_translator (
		.clk                      (clk_clk),                                                              //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                       //                    reset.reset
		.uav_address              (memory_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (memory_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (memory_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (memory_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (memory_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (memory_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (memory_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (memory_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (memory_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (memory_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken                 (memory_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read                  (),                                                                     //              (terminated)
		.av_begintransfer         (),                                                                     //              (terminated)
		.av_beginbursttransfer    (),                                                                     //              (terminated)
		.av_burstcount            (),                                                                     //              (terminated)
		.av_readdatavalid         (1'b0),                                                                 //              (terminated)
		.av_waitrequest           (1'b0),                                                                 //              (terminated)
		.av_writebyteenable       (),                                                                     //              (terminated)
		.av_lock                  (),                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                 //              (terminated)
		.av_debugaccess           (),                                                                     //              (terminated)
		.av_outputenable          (),                                                                     //              (terminated)
		.uav_response             (),                                                                     //              (terminated)
		.av_response              (2'b00),                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ledr_s1_translator (
		.clk                      (clk_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address              (ledr_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ledr_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ledr_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ledr_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ledr_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ledr_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ledr_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ledr_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ledr_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ledr_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ledr_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ledr_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ledr_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ledr_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) uart_0_s1_translator (
		.clk                      (clk_clk),                                                              //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                       //                    reset.reset
		.uav_address              (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (uart_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (uart_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (uart_0_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (uart_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (uart_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (uart_0_s1_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_chipselect            (uart_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_beginbursttransfer    (),                                                                     //              (terminated)
		.av_burstcount            (),                                                                     //              (terminated)
		.av_byteenable            (),                                                                     //              (terminated)
		.av_readdatavalid         (1'b0),                                                                 //              (terminated)
		.av_waitrequest           (1'b0),                                                                 //              (terminated)
		.av_writebyteenable       (),                                                                     //              (terminated)
		.av_lock                  (),                                                                     //              (terminated)
		.av_clken                 (),                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                 //              (terminated)
		.av_debugaccess           (),                                                                     //              (terminated)
		.av_outputenable          (),                                                                     //              (terminated)
		.uav_response             (),                                                                     //              (terminated)
		.av_response              (2'b00),                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                  //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (94),
		.PKT_PROTECTION_L          (92),
		.PKT_BEGIN_BURST           (85),
		.PKT_BURSTWRAP_H           (77),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (80),
		.PKT_BURST_SIZE_L          (78),
		.PKT_BURST_TYPE_H          (82),
		.PKT_BURST_TYPE_L          (81),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (90),
		.PKT_DEST_ID_L             (89),
		.PKT_THREAD_ID_H           (91),
		.PKT_THREAD_ID_L           (91),
		.PKT_CACHE_H               (98),
		.PKT_CACHE_L               (95),
		.PKT_DATA_SIDEBAND_H       (84),
		.PKT_DATA_SIDEBAND_L       (84),
		.PKT_QOS_H                 (86),
		.PKT_QOS_L                 (86),
		.PKT_ADDR_SIDEBAND_H       (83),
		.PKT_ADDR_SIDEBAND_L       (83),
		.PKT_RESPONSE_STATUS_H     (100),
		.PKT_RESPONSE_STATUS_L     (99),
		.ST_DATA_W                 (101),
		.ST_CHANNEL_W              (3),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) rv32i_core_instruction_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                                   //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.av_address              (rv32i_core_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (rv32i_core_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (rv32i_core_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (rv32i_core_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (rv32i_core_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (rv32i_core_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (rv32i_core_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (rv32i_core_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (rv32i_core_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (rv32i_core_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (rv32i_core_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (rv32i_core_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (rv32i_core_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (rv32i_core_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (rv32i_core_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (rv32i_core_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_demux_src0_valid),                                                                 //        rp.valid
		.rp_data                 (rsp_xbar_demux_src0_data),                                                                  //          .data
		.rp_channel              (rsp_xbar_demux_src0_channel),                                                               //          .channel
		.rp_startofpacket        (rsp_xbar_demux_src0_startofpacket),                                                         //          .startofpacket
		.rp_endofpacket          (rsp_xbar_demux_src0_endofpacket),                                                           //          .endofpacket
		.rp_ready                (rsp_xbar_demux_src0_ready),                                                                 //          .ready
		.av_response             (),                                                                                          // (terminated)
		.av_writeresponserequest (1'b0),                                                                                      // (terminated)
		.av_writeresponsevalid   ()                                                                                           // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (94),
		.PKT_PROTECTION_L          (92),
		.PKT_BEGIN_BURST           (85),
		.PKT_BURSTWRAP_H           (77),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (80),
		.PKT_BURST_SIZE_L          (78),
		.PKT_BURST_TYPE_H          (82),
		.PKT_BURST_TYPE_L          (81),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (90),
		.PKT_DEST_ID_L             (89),
		.PKT_THREAD_ID_H           (91),
		.PKT_THREAD_ID_L           (91),
		.PKT_CACHE_H               (98),
		.PKT_CACHE_L               (95),
		.PKT_DATA_SIDEBAND_H       (84),
		.PKT_DATA_SIDEBAND_L       (84),
		.PKT_QOS_H                 (86),
		.PKT_QOS_L                 (86),
		.PKT_ADDR_SIDEBAND_H       (83),
		.PKT_ADDR_SIDEBAND_L       (83),
		.PKT_RESPONSE_STATUS_H     (100),
		.PKT_RESPONSE_STATUS_L     (99),
		.ST_DATA_W                 (101),
		.ST_CHANNEL_W              (3),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) rv32i_core_data_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                            //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.av_address              (rv32i_core_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (rv32i_core_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (rv32i_core_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (rv32i_core_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (rv32i_core_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (rv32i_core_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (rv32i_core_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (rv32i_core_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (rv32i_core_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (rv32i_core_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (rv32i_core_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (rv32i_core_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (rv32i_core_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (rv32i_core_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (rv32i_core_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (rv32i_core_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_001_src_valid),                                                         //        rp.valid
		.rp_data                 (rsp_xbar_mux_001_src_data),                                                          //          .data
		.rp_channel              (rsp_xbar_mux_001_src_channel),                                                       //          .channel
		.rp_startofpacket        (rsp_xbar_mux_001_src_startofpacket),                                                 //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_001_src_endofpacket),                                                   //          .endofpacket
		.rp_ready                (rsp_xbar_mux_001_src_ready),                                                         //          .ready
		.av_response             (),                                                                                   // (terminated)
		.av_writeresponserequest (1'b0),                                                                               // (terminated)
		.av_writeresponsevalid   ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (85),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (90),
		.PKT_DEST_ID_L             (89),
		.PKT_BURSTWRAP_H           (77),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (94),
		.PKT_PROTECTION_L          (92),
		.PKT_RESPONSE_STATUS_H     (100),
		.PKT_RESPONSE_STATUS_L     (99),
		.PKT_BURST_SIZE_H          (80),
		.PKT_BURST_SIZE_L          (78),
		.ST_CHANNEL_W              (3),
		.ST_DATA_W                 (101),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) memory_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (memory_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (memory_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (memory_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (memory_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (memory_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (memory_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (memory_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                       //                .channel
		.rf_sink_ready           (memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (102),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (85),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (90),
		.PKT_DEST_ID_L             (89),
		.PKT_BURSTWRAP_H           (77),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (94),
		.PKT_PROTECTION_L          (92),
		.PKT_RESPONSE_STATUS_H     (100),
		.PKT_RESPONSE_STATUS_L     (99),
		.PKT_BURST_SIZE_H          (80),
		.PKT_BURST_SIZE_L          (78),
		.ST_CHANNEL_W              (3),
		.ST_DATA_W                 (101),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ledr_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (ledr_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ledr_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ledr_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ledr_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ledr_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ledr_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ledr_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ledr_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ledr_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ledr_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ledr_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ledr_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ledr_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ledr_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src1_ready),                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src1_valid),                                                //                .valid
		.cp_data                 (cmd_xbar_demux_001_src1_data),                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src1_startofpacket),                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src1_endofpacket),                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src1_channel),                                              //                .channel
		.rf_sink_ready           (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (102),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (85),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (90),
		.PKT_DEST_ID_L             (89),
		.PKT_BURSTWRAP_H           (77),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (94),
		.PKT_PROTECTION_L          (92),
		.PKT_RESPONSE_STATUS_H     (100),
		.PKT_RESPONSE_STATUS_L     (99),
		.PKT_BURST_SIZE_H          (80),
		.PKT_BURST_SIZE_L          (78),
		.ST_CHANNEL_W              (3),
		.ST_DATA_W                 (101),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) uart_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src2_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src2_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src2_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src2_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src2_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src2_channel),                                                //                .channel
		.rf_sink_ready           (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (102),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	risac_soc_system_addr_router addr_router (
		.sink_ready         (rv32i_core_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (rv32i_core_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (rv32i_core_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (rv32i_core_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (rv32i_core_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                     //       src.ready
		.src_valid          (addr_router_src_valid),                                                                     //          .valid
		.src_data           (addr_router_src_data),                                                                      //          .data
		.src_channel        (addr_router_src_channel),                                                                   //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                             //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                                //          .endofpacket
	);

	risac_soc_system_addr_router_001 addr_router_001 (
		.sink_ready         (rv32i_core_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (rv32i_core_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (rv32i_core_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (rv32i_core_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (rv32i_core_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                          //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                          //          .valid
		.src_data           (addr_router_001_src_data),                                                           //          .data
		.src_channel        (addr_router_001_src_channel),                                                        //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                  //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                     //          .endofpacket
	);

	risac_soc_system_id_router id_router (
		.sink_ready         (memory_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (memory_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (memory_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                  //       src.ready
		.src_valid          (id_router_src_valid),                                                  //          .valid
		.src_data           (id_router_src_data),                                                   //          .data
		.src_channel        (id_router_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                             //          .endofpacket
	);

	risac_soc_system_id_router_001 id_router_001 (
		.sink_ready         (ledr_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ledr_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ledr_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ledr_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ledr_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                            //       src.ready
		.src_valid          (id_router_001_src_valid),                                            //          .valid
		.src_data           (id_router_001_src_data),                                             //          .data
		.src_channel        (id_router_001_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                       //          .endofpacket
	);

	risac_soc_system_id_router_001 id_router_002 (
		.sink_ready         (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                              //       src.ready
		.src_valid          (id_router_002_src_valid),                                              //          .valid
		.src_data           (id_router_002_src_data),                                               //          .data
		.src_channel        (id_router_002_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                         //          .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (clk_clk),                        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

	risac_soc_system_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_src_ready),             //      sink.ready
		.sink_channel       (addr_router_src_channel),           //          .channel
		.sink_data          (addr_router_src_data),              //          .data
		.sink_startofpacket (addr_router_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket)    //          .endofpacket
	);

	risac_soc_system_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_001_src_ready),             //      sink.ready
		.sink_channel       (addr_router_001_src_channel),           //          .channel
		.sink_data          (addr_router_001_src_data),              //          .data
		.sink_startofpacket (addr_router_001_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_001_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_001_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.src2_ready         (cmd_xbar_demux_001_src2_ready),         //      src2.ready
		.src2_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.src2_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.src2_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.src2_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)    //          .endofpacket
	);

	risac_soc_system_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	risac_soc_system_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	risac_soc_system_cmd_xbar_demux rsp_xbar_demux_001 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	risac_soc_system_cmd_xbar_demux rsp_xbar_demux_002 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	risac_soc_system_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

endmodule
