@00000000
93 81 01 00 17 01 02 00 13 01 C1 FF 6F 00 80 0A 
13 01 01 FC 23 24 B1 02 23 26 A1 02 23 22 C1 02 
93 05 00 40 13 06 B0 00 37 05 00 01 23 2C F1 00 
23 2E 11 02 23 2C 51 02 23 2A 61 02 23 28 71 02 
23 20 D1 02 23 2E E1 00 23 2A 01 01 23 28 11 01 
23 26 C1 01 23 24 D1 01 23 22 E1 01 23 20 F1 01 
EF 00 00 0A B7 07 00 03 23 A0 07 00 83 20 C1 03 
83 22 81 03 03 23 41 03 83 23 01 03 03 25 C1 02 
83 25 81 02 03 26 41 02 83 26 01 02 03 27 C1 01 
83 27 81 01 03 28 41 01 83 28 01 01 03 2E C1 00 
83 2E 81 00 03 2F 41 00 83 2F 01 00 13 01 01 04 
73 00 20 30 13 01 01 FF 23 26 11 00 EF 00 C0 06 
93 07 10 00 63 1A F5 02 B3 86 C5 00 37 07 00 01 
63 00 06 02 83 27 47 00 93 D7 07 01 E3 8C 07 FE 
83 C7 05 00 93 85 15 00 23 00 F7 00 E3 94 B6 FE 
13 05 00 00 67 80 00 00 13 05 F0 FF 67 80 00 00 
63 02 06 02 33 87 C5 00 83 27 45 00 93 D7 07 01 
E3 8C 07 FE 83 C7 05 00 93 85 15 00 23 00 F5 00 
E3 14 B7 FE 67 80 00 00 13 01 01 FB 23 26 11 04 
23 24 81 04 23 22 91 04 23 20 21 05 23 2E 31 03 
23 2C 41 03 23 2A 51 03 23 28 61 03 23 26 71 03 
23 24 81 03 23 22 91 03 23 20 A1 03 B7 07 00 02 
13 07 00 05 23 80 E7 00 93 07 00 01 73 90 57 30 
93 07 00 08 73 A0 47 30 13 07 40 41 F3 27 50 30 
03 2A 07 00 83 29 47 00 03 29 87 00 83 24 C7 00 
03 44 07 01 13 D7 87 00 13 77 F7 0F 93 D5 87 01 
13 58 47 00 93 06 01 02 13 77 F7 00 33 88 06 01 
13 D6 07 01 B3 86 E6 00 13 D5 C7 01 13 07 01 02 
93 F5 F5 00 23 26 41 01 23 28 31 01 23 2A 21 01 
23 2C 91 00 23 0E 81 00 33 05 A7 00 B3 05 B7 00 
13 76 F6 0F 93 F7 F7 0F 03 47 C8 FE 03 C3 C6 FE 
83 C8 C5 FE 83 46 C5 FE 13 08 01 02 13 D5 47 00 
93 55 46 00 B3 05 B8 00 33 05 A8 00 37 0D FF FF 
03 48 C5 FE 13 0D FD 0F 03 C5 C5 FE 93 F7 F7 00 
93 05 01 02 13 76 F6 00 13 13 83 00 93 98 88 00 
33 77 A7 01 B3 87 F5 00 B3 F6 A6 01 33 86 C5 00 
B7 0C 01 FF 83 C5 C7 FE 03 46 C6 FE B3 67 67 00 
93 8C FC FF 33 E7 16 01 13 18 08 01 93 16 05 01 
B3 F7 97 01 33 77 97 01 37 0C 00 01 B3 E7 07 01 
13 0C FC FF 33 67 D7 00 93 95 85 01 93 16 86 01 
B3 F7 87 01 33 77 87 01 B3 E7 B7 00 33 67 D7 00 
13 06 20 00 93 05 C0 40 37 05 00 01 23 24 F1 00 
23 22 E1 00 EF F0 DF E5 13 06 80 00 93 05 41 00 
37 05 00 01 EF F0 DF E4 13 06 10 00 93 05 00 41 
37 05 00 01 EF F0 DF E3 B7 07 00 03 13 06 00 50 
93 06 00 00 23 A4 C7 00 23 A6 D7 00 93 0B 00 00 
93 D7 8B 00 93 F7 F7 0F 93 D5 8B 01 13 D8 47 00 
13 07 01 02 93 F7 F7 00 33 08 07 01 93 D6 0B 01 
33 07 F7 00 13 D5 CB 01 93 07 01 02 93 F5 F5 00 
23 26 41 01 23 28 31 01 23 2A 21 01 23 2C 91 00 
23 0E 81 00 13 F6 FB 0F 33 85 A7 00 B3 85 B7 00 
93 F6 F6 0F 13 03 01 02 83 47 C8 FE 83 48 C7 FE 
03 C8 C5 FE 03 47 C5 FE 93 D5 46 00 13 55 46 00 
33 05 A3 00 B3 05 B3 00 03 45 C5 FE 83 C5 C5 FE 
13 76 F6 00 93 F6 F6 00 93 98 88 00 33 06 C3 00 
13 18 88 00 B3 06 D3 00 B3 F7 A7 01 33 77 A7 01 
B3 E7 17 01 33 67 07 01 03 46 C6 FE 83 C6 C6 FE 
13 15 05 01 93 95 05 01 B3 F7 97 01 33 77 97 01 
B3 E7 A7 00 33 67 B7 00 93 96 86 01 13 16 86 01 
B3 F7 87 01 33 77 87 01 B3 E7 C7 00 33 67 D7 00 
13 06 20 00 93 05 C0 40 37 05 00 01 23 22 E1 00 
23 24 F1 00 EF F0 DF D2 13 06 80 00 93 05 41 00 
37 05 00 01 EF F0 DF D1 13 06 10 00 93 05 00 41 
37 05 00 01 EF F0 DF D0 93 8B 1B 00 6F F0 5F EE 
@00000400
49 54 53 20 41 20 54 52 41 50 00 00 30 78 00 00 
0A 00 00 00 30 31 32 33 34 35 36 37 38 39 61 62 
63 64 65 66 00 00 00 00 
