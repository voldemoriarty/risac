library verilog;
use verilog.vl_types.all;
entity risac_soc_tb is
end risac_soc_tb;
