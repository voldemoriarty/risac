@00000000
17 11 00 00 13 01 01 00 6F 00 40 00 13 01 01 FF 
23 26 11 00 EF 00 40 00 37 07 00 02 93 06 50 05 
93 07 40 04 23 00 D7 00 93 86 37 01 37 07 00 01 
03 C6 07 00 93 87 17 00 23 00 C7 00 E3 9A D7 FE 
6F 00 00 00 
@00000044
57 65 6C 63 6F 6D 65 20 44 72 20 41 77 61 69 73 
0D 0A 00 00 
