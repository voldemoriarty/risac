@00000000
17 11 00 00 13 01 01 00 6F 00 40 00 13 01 01 FF 
23 26 11 00 EF 00 40 00 13 07 50 05 93 06 00 05 
B7 07 00 02 23 80 E7 00 13 86 36 01 37 07 00 01 
83 27 47 00 93 D7 07 01 E3 8C 07 FE 83 C7 06 00 
93 86 16 00 23 00 F7 00 E3 94 C6 FE 6F 00 00 00 
@00000050
57 65 6C 63 6F 6D 65 20 44 72 20 41 77 61 69 73 
0D 0A 00 00 
