@00000000
93 81 01 00 17 01 02 00 13 01 C1 FF 6F 00 00 0A 
13 01 01 FC 23 24 B1 02 23 26 A1 02 23 22 C1 02 
93 05 C0 28 13 06 B0 00 37 05 00 01 23 2E 11 02 
23 2C 51 02 23 2A 61 02 23 28 71 02 23 20 D1 02 
23 2E E1 00 23 2C F1 00 23 2A 01 01 23 28 11 01 
23 26 C1 01 23 24 D1 01 23 22 E1 01 23 20 F1 01 
EF 00 80 05 83 20 C1 03 83 22 81 03 03 23 41 03 
83 23 01 03 03 25 C1 02 83 25 81 02 03 26 41 02 
83 26 01 02 03 27 C1 01 83 27 81 01 03 28 41 01 
83 28 01 01 03 2E C1 00 83 2E 81 00 03 2F 41 00 
83 2F 01 00 13 01 01 04 73 00 20 30 13 01 01 FF 
23 26 11 00 EF 00 00 06 93 07 00 00 63 94 C7 00 
67 80 00 00 03 27 45 00 13 57 07 01 E3 0C 07 FE 
33 87 F5 00 03 47 07 00 93 87 17 00 23 00 E5 00 
6F F0 DF FD 93 07 10 00 63 12 F5 02 13 01 01 FF 
37 05 00 01 23 26 11 00 EF F0 1F FC 83 20 C1 00 
13 05 00 00 13 01 01 01 67 80 00 00 13 05 F0 FF 
67 80 00 00 13 01 01 FD 23 26 11 02 B7 07 00 02 
13 07 00 05 23 80 E7 00 93 07 00 01 73 90 57 30 
93 07 00 08 73 A0 47 30 13 07 C0 29 83 46 07 01 
F3 27 50 30 83 2E 07 00 03 2E 47 00 03 23 87 00 
83 28 C7 00 13 D7 87 00 13 77 F7 0F 23 0E D1 00 
93 D5 87 01 13 58 47 00 93 06 01 02 13 77 F7 00 
33 88 06 01 13 D6 07 01 B3 86 E6 00 13 D5 C7 01 
13 07 01 02 93 F5 F5 00 23 26 D1 01 23 28 C1 01 
23 2A 61 00 23 2C 11 01 33 05 A7 00 B3 05 B7 00 
13 76 F6 0F 93 F7 F7 0F 03 47 C8 FE 03 CE C6 FE 
03 C3 C5 FE 83 46 C5 FE 93 05 01 02 13 D8 47 00 
13 55 46 00 33 88 05 01 33 85 A5 00 B7 05 FF FF 
83 48 C8 FE 93 85 F5 0F 03 48 C5 FE 93 F7 F7 00 
13 05 01 02 13 1E 8E 00 33 77 B7 00 B3 F6 B6 00 
B3 07 F5 00 13 76 F6 00 B7 05 01 FF 13 13 83 00 
93 85 F5 FF 33 06 C5 00 03 C5 C7 FE B3 67 C7 01 
93 98 08 01 33 E7 66 00 03 46 C6 FE B3 F7 B7 00 
B7 06 00 01 93 86 F6 FF 13 18 08 01 B3 E7 17 01 
33 77 B7 00 33 67 07 01 93 15 85 01 B3 F7 D7 00 
B3 E7 B7 00 33 77 D7 00 13 16 86 01 33 67 C7 00 
93 05 80 29 13 06 20 00 37 05 00 01 23 22 E1 00 
23 24 F1 00 EF F0 5F E5 13 06 80 00 93 05 41 00 
37 05 00 01 EF F0 5F E4 B7 07 00 03 13 07 00 50 
23 A4 E7 00 23 A6 07 00 6F 00 00 00 
@0000028C
49 54 53 20 41 20 54 52 41 50 00 00 30 78 00 00 
30 31 32 33 34 35 36 37 38 39 61 62 63 64 65 66 
00 00 00 00 
