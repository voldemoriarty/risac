@00000000
17 11 00 00 13 01 01 00 6F 00 C0 02 63 52 C0 02 
33 87 C5 00 83 27 45 00 93 D7 07 01 E3 8C 07 FE 
83 C7 05 00 93 85 15 00 23 00 F5 00 E3 94 E5 FE 
67 80 00 00 13 01 01 FF 23 26 11 00 EF 00 40 00 
B7 07 00 02 13 07 00 05 23 80 E7 00 B7 77 6C 6F 
13 01 01 FF 93 87 57 C6 23 24 F1 00 B7 17 00 00 
93 87 D7 A0 23 16 F1 00 23 07 01 00 93 06 81 00 
13 06 F1 00 37 07 00 01 83 27 47 00 93 D7 07 01 
E3 8C 07 FE 83 C7 06 00 93 86 16 00 23 00 F7 00 
E3 94 C6 FE 6F 00 00 00 
