@00000000
17 11 00 00 13 01 01 00 6F 00 C0 02 63 52 C0 02 
33 87 C5 00 83 27 45 00 93 D7 07 01 E3 8C 07 FE 
83 C7 05 00 93 85 15 00 23 00 F5 00 E3 94 E5 FE 
67 80 00 00 13 01 01 FF 23 26 11 00 EF 00 40 00 
13 07 50 05 B7 07 00 02 23 80 E7 00 93 05 C0 07 
13 06 C0 08 37 07 00 01 93 86 05 00 83 27 47 00 
93 D7 07 01 E3 8C 07 FE 83 C7 06 00 93 86 16 00 
23 00 F7 00 E3 94 C6 FE 6F F0 1F FE 
@0000007C
48 65 6C 6C 6F 2C 20 57 6F 72 6C 64 21 0D 0A 00 
