@00000000
B7 17 00 00 83 A7 07 00 13 81 07 00 6F 00 40 00 
13 01 01 FF 23 26 11 00 EF 00 40 00 B7 07 01 00 
13 07 80 04 23 80 E7 00 13 07 50 06 23 80 E7 00 
13 07 C0 06 23 80 E7 00 23 80 E7 00 93 06 F0 06 
23 80 D7 00 13 06 C0 02 23 80 C7 00 13 06 00 02 
23 80 C7 00 13 06 70 05 23 80 C7 00 23 80 D7 00 
93 06 20 07 23 80 D7 00 23 80 E7 00 13 07 40 06 
23 80 E7 00 13 07 10 02 23 80 E7 00 13 07 A0 00 
23 80 E7 00 37 87 01 00 13 01 01 FF 23 80 07 00 
93 06 00 00 13 07 F7 69 23 26 01 00 83 27 C1 00 
63 6C F7 00 83 27 C1 00 93 87 17 00 23 26 F1 00 
83 27 C1 00 E3 78 F7 FE 23 24 01 00 83 27 81 00 
63 6C F7 00 83 27 81 00 93 87 17 00 23 24 F1 00 
83 27 81 00 E3 78 F7 FE 23 24 D0 00 93 86 16 00 
6F F0 9F FB 
